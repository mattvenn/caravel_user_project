magic
tech sky130A
magscale 1 2
timestamp 1619619845
<< obsli1 >>
rect 69904 94959 514080 608881
<< obsm1 >>
rect 566 1640 582820 702704
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 572 703464 8030 703520
rect 8254 703464 24222 703520
rect 24446 703464 40414 703520
rect 40638 703464 56698 703520
rect 56922 703464 72890 703520
rect 73114 703464 89082 703520
rect 89306 703464 105366 703520
rect 105590 703464 121558 703520
rect 121782 703464 137750 703520
rect 137974 703464 154034 703520
rect 154258 703464 170226 703520
rect 170450 703464 186418 703520
rect 186642 703464 202702 703520
rect 202926 703464 218894 703520
rect 219118 703464 235086 703520
rect 235310 703464 251370 703520
rect 251594 703464 267562 703520
rect 267786 703464 283754 703520
rect 283978 703464 300038 703520
rect 300262 703464 316230 703520
rect 316454 703464 332422 703520
rect 332646 703464 348706 703520
rect 348930 703464 364898 703520
rect 365122 703464 381090 703520
rect 381314 703464 397374 703520
rect 397598 703464 413566 703520
rect 413790 703464 429758 703520
rect 429982 703464 446042 703520
rect 446266 703464 462234 703520
rect 462458 703464 478426 703520
rect 478650 703464 494710 703520
rect 494934 703464 510902 703520
rect 511126 703464 527094 703520
rect 527318 703464 543378 703520
rect 543602 703464 559570 703520
rect 559794 703464 575762 703520
rect 575986 703464 580410 703520
rect 572 536 580410 703464
rect 710 480 1590 536
rect 1814 480 2786 536
rect 3010 480 3982 536
rect 4206 480 5178 536
rect 5402 480 6374 536
rect 6598 480 7570 536
rect 7794 480 8766 536
rect 8990 480 9962 536
rect 10186 480 11158 536
rect 11382 480 12354 536
rect 12578 480 13550 536
rect 13774 480 14746 536
rect 14970 480 15942 536
rect 16166 480 17138 536
rect 17362 480 18242 536
rect 18466 480 19438 536
rect 19662 480 20634 536
rect 20858 480 21830 536
rect 22054 480 23026 536
rect 23250 480 24222 536
rect 24446 480 25418 536
rect 25642 480 26614 536
rect 26838 480 27810 536
rect 28034 480 29006 536
rect 29230 480 30202 536
rect 30426 480 31398 536
rect 31622 480 32594 536
rect 32818 480 33790 536
rect 34014 480 34894 536
rect 35118 480 36090 536
rect 36314 480 37286 536
rect 37510 480 38482 536
rect 38706 480 39678 536
rect 39902 480 40874 536
rect 41098 480 42070 536
rect 42294 480 43266 536
rect 43490 480 44462 536
rect 44686 480 45658 536
rect 45882 480 46854 536
rect 47078 480 48050 536
rect 48274 480 49246 536
rect 49470 480 50442 536
rect 50666 480 51546 536
rect 51770 480 52742 536
rect 52966 480 53938 536
rect 54162 480 55134 536
rect 55358 480 56330 536
rect 56554 480 57526 536
rect 57750 480 58722 536
rect 58946 480 59918 536
rect 60142 480 61114 536
rect 61338 480 62310 536
rect 62534 480 63506 536
rect 63730 480 64702 536
rect 64926 480 65898 536
rect 66122 480 67094 536
rect 67318 480 68198 536
rect 68422 480 69394 536
rect 69618 480 70590 536
rect 70814 480 71786 536
rect 72010 480 72982 536
rect 73206 480 74178 536
rect 74402 480 75374 536
rect 75598 480 76570 536
rect 76794 480 77766 536
rect 77990 480 78962 536
rect 79186 480 80158 536
rect 80382 480 81354 536
rect 81578 480 82550 536
rect 82774 480 83746 536
rect 83970 480 84850 536
rect 85074 480 86046 536
rect 86270 480 87242 536
rect 87466 480 88438 536
rect 88662 480 89634 536
rect 89858 480 90830 536
rect 91054 480 92026 536
rect 92250 480 93222 536
rect 93446 480 94418 536
rect 94642 480 95614 536
rect 95838 480 96810 536
rect 97034 480 98006 536
rect 98230 480 99202 536
rect 99426 480 100398 536
rect 100622 480 101502 536
rect 101726 480 102698 536
rect 102922 480 103894 536
rect 104118 480 105090 536
rect 105314 480 106286 536
rect 106510 480 107482 536
rect 107706 480 108678 536
rect 108902 480 109874 536
rect 110098 480 111070 536
rect 111294 480 112266 536
rect 112490 480 113462 536
rect 113686 480 114658 536
rect 114882 480 115854 536
rect 116078 480 117050 536
rect 117274 480 118154 536
rect 118378 480 119350 536
rect 119574 480 120546 536
rect 120770 480 121742 536
rect 121966 480 122938 536
rect 123162 480 124134 536
rect 124358 480 125330 536
rect 125554 480 126526 536
rect 126750 480 127722 536
rect 127946 480 128918 536
rect 129142 480 130114 536
rect 130338 480 131310 536
rect 131534 480 132506 536
rect 132730 480 133702 536
rect 133926 480 134806 536
rect 135030 480 136002 536
rect 136226 480 137198 536
rect 137422 480 138394 536
rect 138618 480 139590 536
rect 139814 480 140786 536
rect 141010 480 141982 536
rect 142206 480 143178 536
rect 143402 480 144374 536
rect 144598 480 145570 536
rect 145794 480 146766 536
rect 146990 480 147962 536
rect 148186 480 149158 536
rect 149382 480 150354 536
rect 150578 480 151458 536
rect 151682 480 152654 536
rect 152878 480 153850 536
rect 154074 480 155046 536
rect 155270 480 156242 536
rect 156466 480 157438 536
rect 157662 480 158634 536
rect 158858 480 159830 536
rect 160054 480 161026 536
rect 161250 480 162222 536
rect 162446 480 163418 536
rect 163642 480 164614 536
rect 164838 480 165810 536
rect 166034 480 167006 536
rect 167230 480 168110 536
rect 168334 480 169306 536
rect 169530 480 170502 536
rect 170726 480 171698 536
rect 171922 480 172894 536
rect 173118 480 174090 536
rect 174314 480 175286 536
rect 175510 480 176482 536
rect 176706 480 177678 536
rect 177902 480 178874 536
rect 179098 480 180070 536
rect 180294 480 181266 536
rect 181490 480 182462 536
rect 182686 480 183658 536
rect 183882 480 184762 536
rect 184986 480 185958 536
rect 186182 480 187154 536
rect 187378 480 188350 536
rect 188574 480 189546 536
rect 189770 480 190742 536
rect 190966 480 191938 536
rect 192162 480 193134 536
rect 193358 480 194330 536
rect 194554 480 195526 536
rect 195750 480 196722 536
rect 196946 480 197918 536
rect 198142 480 199114 536
rect 199338 480 200310 536
rect 200534 480 201414 536
rect 201638 480 202610 536
rect 202834 480 203806 536
rect 204030 480 205002 536
rect 205226 480 206198 536
rect 206422 480 207394 536
rect 207618 480 208590 536
rect 208814 480 209786 536
rect 210010 480 210982 536
rect 211206 480 212178 536
rect 212402 480 213374 536
rect 213598 480 214570 536
rect 214794 480 215766 536
rect 215990 480 216962 536
rect 217186 480 218066 536
rect 218290 480 219262 536
rect 219486 480 220458 536
rect 220682 480 221654 536
rect 221878 480 222850 536
rect 223074 480 224046 536
rect 224270 480 225242 536
rect 225466 480 226438 536
rect 226662 480 227634 536
rect 227858 480 228830 536
rect 229054 480 230026 536
rect 230250 480 231222 536
rect 231446 480 232418 536
rect 232642 480 233614 536
rect 233838 480 234718 536
rect 234942 480 235914 536
rect 236138 480 237110 536
rect 237334 480 238306 536
rect 238530 480 239502 536
rect 239726 480 240698 536
rect 240922 480 241894 536
rect 242118 480 243090 536
rect 243314 480 244286 536
rect 244510 480 245482 536
rect 245706 480 246678 536
rect 246902 480 247874 536
rect 248098 480 249070 536
rect 249294 480 250266 536
rect 250490 480 251370 536
rect 251594 480 252566 536
rect 252790 480 253762 536
rect 253986 480 254958 536
rect 255182 480 256154 536
rect 256378 480 257350 536
rect 257574 480 258546 536
rect 258770 480 259742 536
rect 259966 480 260938 536
rect 261162 480 262134 536
rect 262358 480 263330 536
rect 263554 480 264526 536
rect 264750 480 265722 536
rect 265946 480 266918 536
rect 267142 480 268022 536
rect 268246 480 269218 536
rect 269442 480 270414 536
rect 270638 480 271610 536
rect 271834 480 272806 536
rect 273030 480 274002 536
rect 274226 480 275198 536
rect 275422 480 276394 536
rect 276618 480 277590 536
rect 277814 480 278786 536
rect 279010 480 279982 536
rect 280206 480 281178 536
rect 281402 480 282374 536
rect 282598 480 283570 536
rect 283794 480 284674 536
rect 284898 480 285870 536
rect 286094 480 287066 536
rect 287290 480 288262 536
rect 288486 480 289458 536
rect 289682 480 290654 536
rect 290878 480 291850 536
rect 292074 480 293046 536
rect 293270 480 294242 536
rect 294466 480 295438 536
rect 295662 480 296634 536
rect 296858 480 297830 536
rect 298054 480 299026 536
rect 299250 480 300222 536
rect 300446 480 301326 536
rect 301550 480 302522 536
rect 302746 480 303718 536
rect 303942 480 304914 536
rect 305138 480 306110 536
rect 306334 480 307306 536
rect 307530 480 308502 536
rect 308726 480 309698 536
rect 309922 480 310894 536
rect 311118 480 312090 536
rect 312314 480 313286 536
rect 313510 480 314482 536
rect 314706 480 315678 536
rect 315902 480 316874 536
rect 317098 480 317978 536
rect 318202 480 319174 536
rect 319398 480 320370 536
rect 320594 480 321566 536
rect 321790 480 322762 536
rect 322986 480 323958 536
rect 324182 480 325154 536
rect 325378 480 326350 536
rect 326574 480 327546 536
rect 327770 480 328742 536
rect 328966 480 329938 536
rect 330162 480 331134 536
rect 331358 480 332330 536
rect 332554 480 333526 536
rect 333750 480 334630 536
rect 334854 480 335826 536
rect 336050 480 337022 536
rect 337246 480 338218 536
rect 338442 480 339414 536
rect 339638 480 340610 536
rect 340834 480 341806 536
rect 342030 480 343002 536
rect 343226 480 344198 536
rect 344422 480 345394 536
rect 345618 480 346590 536
rect 346814 480 347786 536
rect 348010 480 348982 536
rect 349206 480 350178 536
rect 350402 480 351282 536
rect 351506 480 352478 536
rect 352702 480 353674 536
rect 353898 480 354870 536
rect 355094 480 356066 536
rect 356290 480 357262 536
rect 357486 480 358458 536
rect 358682 480 359654 536
rect 359878 480 360850 536
rect 361074 480 362046 536
rect 362270 480 363242 536
rect 363466 480 364438 536
rect 364662 480 365634 536
rect 365858 480 366830 536
rect 367054 480 367934 536
rect 368158 480 369130 536
rect 369354 480 370326 536
rect 370550 480 371522 536
rect 371746 480 372718 536
rect 372942 480 373914 536
rect 374138 480 375110 536
rect 375334 480 376306 536
rect 376530 480 377502 536
rect 377726 480 378698 536
rect 378922 480 379894 536
rect 380118 480 381090 536
rect 381314 480 382286 536
rect 382510 480 383482 536
rect 383706 480 384586 536
rect 384810 480 385782 536
rect 386006 480 386978 536
rect 387202 480 388174 536
rect 388398 480 389370 536
rect 389594 480 390566 536
rect 390790 480 391762 536
rect 391986 480 392958 536
rect 393182 480 394154 536
rect 394378 480 395350 536
rect 395574 480 396546 536
rect 396770 480 397742 536
rect 397966 480 398938 536
rect 399162 480 400134 536
rect 400358 480 401238 536
rect 401462 480 402434 536
rect 402658 480 403630 536
rect 403854 480 404826 536
rect 405050 480 406022 536
rect 406246 480 407218 536
rect 407442 480 408414 536
rect 408638 480 409610 536
rect 409834 480 410806 536
rect 411030 480 412002 536
rect 412226 480 413198 536
rect 413422 480 414394 536
rect 414618 480 415590 536
rect 415814 480 416786 536
rect 417010 480 417890 536
rect 418114 480 419086 536
rect 419310 480 420282 536
rect 420506 480 421478 536
rect 421702 480 422674 536
rect 422898 480 423870 536
rect 424094 480 425066 536
rect 425290 480 426262 536
rect 426486 480 427458 536
rect 427682 480 428654 536
rect 428878 480 429850 536
rect 430074 480 431046 536
rect 431270 480 432242 536
rect 432466 480 433438 536
rect 433662 480 434542 536
rect 434766 480 435738 536
rect 435962 480 436934 536
rect 437158 480 438130 536
rect 438354 480 439326 536
rect 439550 480 440522 536
rect 440746 480 441718 536
rect 441942 480 442914 536
rect 443138 480 444110 536
rect 444334 480 445306 536
rect 445530 480 446502 536
rect 446726 480 447698 536
rect 447922 480 448894 536
rect 449118 480 450090 536
rect 450314 480 451194 536
rect 451418 480 452390 536
rect 452614 480 453586 536
rect 453810 480 454782 536
rect 455006 480 455978 536
rect 456202 480 457174 536
rect 457398 480 458370 536
rect 458594 480 459566 536
rect 459790 480 460762 536
rect 460986 480 461958 536
rect 462182 480 463154 536
rect 463378 480 464350 536
rect 464574 480 465546 536
rect 465770 480 466742 536
rect 466966 480 467846 536
rect 468070 480 469042 536
rect 469266 480 470238 536
rect 470462 480 471434 536
rect 471658 480 472630 536
rect 472854 480 473826 536
rect 474050 480 475022 536
rect 475246 480 476218 536
rect 476442 480 477414 536
rect 477638 480 478610 536
rect 478834 480 479806 536
rect 480030 480 481002 536
rect 481226 480 482198 536
rect 482422 480 483394 536
rect 483618 480 484498 536
rect 484722 480 485694 536
rect 485918 480 486890 536
rect 487114 480 488086 536
rect 488310 480 489282 536
rect 489506 480 490478 536
rect 490702 480 491674 536
rect 491898 480 492870 536
rect 493094 480 494066 536
rect 494290 480 495262 536
rect 495486 480 496458 536
rect 496682 480 497654 536
rect 497878 480 498850 536
rect 499074 480 500046 536
rect 500270 480 501150 536
rect 501374 480 502346 536
rect 502570 480 503542 536
rect 503766 480 504738 536
rect 504962 480 505934 536
rect 506158 480 507130 536
rect 507354 480 508326 536
rect 508550 480 509522 536
rect 509746 480 510718 536
rect 510942 480 511914 536
rect 512138 480 513110 536
rect 513334 480 514306 536
rect 514530 480 515502 536
rect 515726 480 516698 536
rect 516922 480 517802 536
rect 518026 480 518998 536
rect 519222 480 520194 536
rect 520418 480 521390 536
rect 521614 480 522586 536
rect 522810 480 523782 536
rect 524006 480 524978 536
rect 525202 480 526174 536
rect 526398 480 527370 536
rect 527594 480 528566 536
rect 528790 480 529762 536
rect 529986 480 530958 536
rect 531182 480 532154 536
rect 532378 480 533350 536
rect 533574 480 534454 536
rect 534678 480 535650 536
rect 535874 480 536846 536
rect 537070 480 538042 536
rect 538266 480 539238 536
rect 539462 480 540434 536
rect 540658 480 541630 536
rect 541854 480 542826 536
rect 543050 480 544022 536
rect 544246 480 545218 536
rect 545442 480 546414 536
rect 546638 480 547610 536
rect 547834 480 548806 536
rect 549030 480 550002 536
rect 550226 480 551106 536
rect 551330 480 552302 536
rect 552526 480 553498 536
rect 553722 480 554694 536
rect 554918 480 555890 536
rect 556114 480 557086 536
rect 557310 480 558282 536
rect 558506 480 559478 536
rect 559702 480 560674 536
rect 560898 480 561870 536
rect 562094 480 563066 536
rect 563290 480 564262 536
rect 564486 480 565458 536
rect 565682 480 566654 536
rect 566878 480 567758 536
rect 567982 480 568954 536
rect 569178 480 570150 536
rect 570374 480 571346 536
rect 571570 480 572542 536
rect 572766 480 573738 536
rect 573962 480 574934 536
rect 575158 480 576130 536
rect 576354 480 577326 536
rect 577550 480 578522 536
rect 578746 480 579718 536
rect 579942 480 580410 536
<< metal3 >>
rect 583520 697900 584960 698140
rect -960 696268 480 696508
rect 583520 686204 584960 686444
rect -960 681308 480 681548
rect 583520 674508 584960 674748
rect -960 666348 480 666588
rect 583520 662676 584960 662916
rect -960 651388 480 651628
rect 583520 650980 584960 651220
rect 583520 639284 584960 639524
rect -960 636428 480 636668
rect 583520 627588 584960 627828
rect -960 621468 480 621708
rect 583520 615756 584960 615996
rect -960 606508 480 606748
rect 583520 604060 584960 604300
rect 583520 592364 584960 592604
rect -960 591412 480 591652
rect 583520 580668 584960 580908
rect -960 576452 480 576692
rect 583520 568836 584960 569076
rect -960 561492 480 561732
rect 583520 557140 584960 557380
rect -960 546532 480 546772
rect 583520 545444 584960 545684
rect 583520 533748 584960 533988
rect -960 531572 480 531812
rect 583520 521916 584960 522156
rect -960 516612 480 516852
rect 583520 510220 584960 510460
rect -960 501652 480 501892
rect 583520 498524 584960 498764
rect -960 486692 480 486932
rect 583520 486692 584960 486932
rect 583520 474996 584960 475236
rect -960 471596 480 471836
rect 583520 463300 584960 463540
rect -960 456636 480 456876
rect 583520 451604 584960 451844
rect -960 441676 480 441916
rect 583520 439772 584960 440012
rect 583520 428076 584960 428316
rect -960 426716 480 426956
rect 583520 416380 584960 416620
rect -960 411756 480 411996
rect 583520 404684 584960 404924
rect -960 396796 480 397036
rect 583520 392852 584960 393092
rect -960 381836 480 382076
rect 583520 381156 584960 381396
rect 583520 369460 584960 369700
rect -960 366876 480 367116
rect 583520 357764 584960 358004
rect -960 351780 480 352020
rect 583520 345932 584960 346172
rect -960 336820 480 337060
rect 583520 334236 584960 334476
rect 583520 322540 584960 322780
rect -960 321860 480 322100
rect 583520 310708 584960 310948
rect -960 306900 480 307140
rect 583520 299012 584960 299252
rect -960 291940 480 292180
rect 583520 287316 584960 287556
rect -960 276980 480 277220
rect 583520 275620 584960 275860
rect 583520 263788 584960 264028
rect -960 262020 480 262260
rect 583520 252092 584960 252332
rect -960 247060 480 247300
rect 583520 240396 584960 240636
rect -960 231964 480 232204
rect 583520 228700 584960 228940
rect -960 217004 480 217244
rect 583520 216868 584960 217108
rect 583520 205172 584960 205412
rect -960 202044 480 202284
rect 583520 193476 584960 193716
rect -960 187084 480 187324
rect 583520 181780 584960 182020
rect -960 172124 480 172364
rect 583520 169948 584960 170188
rect 583520 158252 584960 158492
rect -960 157164 480 157404
rect 583520 146556 584960 146796
rect -960 142204 480 142444
rect 583520 134724 584960 134964
rect -960 127244 480 127484
rect 583520 123028 584960 123268
rect -960 112148 480 112388
rect 583520 111332 584960 111572
rect 583520 99636 584960 99876
rect -960 97188 480 97428
rect 583520 87804 584960 88044
rect -960 82228 480 82468
rect 583520 76108 584960 76348
rect -960 67268 480 67508
rect 583520 64412 584960 64652
rect 583520 52716 584960 52956
rect -960 52308 480 52548
rect 583520 40884 584960 41124
rect -960 37348 480 37588
rect 583520 29188 584960 29428
rect -960 22388 480 22628
rect 583520 17492 584960 17732
rect -960 7428 480 7668
rect 583520 5796 584960 6036
<< obsm3 >>
rect 480 698220 583520 702541
rect 480 697820 583440 698220
rect 480 696588 583520 697820
rect 560 696188 583520 696588
rect 480 686524 583520 696188
rect 480 686124 583440 686524
rect 480 681628 583520 686124
rect 560 681228 583520 681628
rect 480 674828 583520 681228
rect 480 674428 583440 674828
rect 480 666668 583520 674428
rect 560 666268 583520 666668
rect 480 662996 583520 666268
rect 480 662596 583440 662996
rect 480 651708 583520 662596
rect 560 651308 583520 651708
rect 480 651300 583520 651308
rect 480 650900 583440 651300
rect 480 639604 583520 650900
rect 480 639204 583440 639604
rect 480 636748 583520 639204
rect 560 636348 583520 636748
rect 480 627908 583520 636348
rect 480 627508 583440 627908
rect 480 621788 583520 627508
rect 560 621388 583520 621788
rect 480 616076 583520 621388
rect 480 615676 583440 616076
rect 480 606828 583520 615676
rect 560 606428 583520 606828
rect 480 604380 583520 606428
rect 480 603980 583440 604380
rect 480 592684 583520 603980
rect 480 592284 583440 592684
rect 480 591732 583520 592284
rect 560 591332 583520 591732
rect 480 580988 583520 591332
rect 480 580588 583440 580988
rect 480 576772 583520 580588
rect 560 576372 583520 576772
rect 480 569156 583520 576372
rect 480 568756 583440 569156
rect 480 561812 583520 568756
rect 560 561412 583520 561812
rect 480 557460 583520 561412
rect 480 557060 583440 557460
rect 480 546852 583520 557060
rect 560 546452 583520 546852
rect 480 545764 583520 546452
rect 480 545364 583440 545764
rect 480 534068 583520 545364
rect 480 533668 583440 534068
rect 480 531892 583520 533668
rect 560 531492 583520 531892
rect 480 522236 583520 531492
rect 480 521836 583440 522236
rect 480 516932 583520 521836
rect 560 516532 583520 516932
rect 480 510540 583520 516532
rect 480 510140 583440 510540
rect 480 501972 583520 510140
rect 560 501572 583520 501972
rect 480 498844 583520 501572
rect 480 498444 583440 498844
rect 480 487012 583520 498444
rect 560 486612 583440 487012
rect 480 475316 583520 486612
rect 480 474916 583440 475316
rect 480 471916 583520 474916
rect 560 471516 583520 471916
rect 480 463620 583520 471516
rect 480 463220 583440 463620
rect 480 456956 583520 463220
rect 560 456556 583520 456956
rect 480 451924 583520 456556
rect 480 451524 583440 451924
rect 480 441996 583520 451524
rect 560 441596 583520 441996
rect 480 440092 583520 441596
rect 480 439692 583440 440092
rect 480 428396 583520 439692
rect 480 427996 583440 428396
rect 480 427036 583520 427996
rect 560 426636 583520 427036
rect 480 416700 583520 426636
rect 480 416300 583440 416700
rect 480 412076 583520 416300
rect 560 411676 583520 412076
rect 480 405004 583520 411676
rect 480 404604 583440 405004
rect 480 397116 583520 404604
rect 560 396716 583520 397116
rect 480 393172 583520 396716
rect 480 392772 583440 393172
rect 480 382156 583520 392772
rect 560 381756 583520 382156
rect 480 381476 583520 381756
rect 480 381076 583440 381476
rect 480 369780 583520 381076
rect 480 369380 583440 369780
rect 480 367196 583520 369380
rect 560 366796 583520 367196
rect 480 358084 583520 366796
rect 480 357684 583440 358084
rect 480 352100 583520 357684
rect 560 351700 583520 352100
rect 480 346252 583520 351700
rect 480 345852 583440 346252
rect 480 337140 583520 345852
rect 560 336740 583520 337140
rect 480 334556 583520 336740
rect 480 334156 583440 334556
rect 480 322860 583520 334156
rect 480 322460 583440 322860
rect 480 322180 583520 322460
rect 560 321780 583520 322180
rect 480 311028 583520 321780
rect 480 310628 583440 311028
rect 480 307220 583520 310628
rect 560 306820 583520 307220
rect 480 299332 583520 306820
rect 480 298932 583440 299332
rect 480 292260 583520 298932
rect 560 291860 583520 292260
rect 480 287636 583520 291860
rect 480 287236 583440 287636
rect 480 277300 583520 287236
rect 560 276900 583520 277300
rect 480 275940 583520 276900
rect 480 275540 583440 275940
rect 480 264108 583520 275540
rect 480 263708 583440 264108
rect 480 262340 583520 263708
rect 560 261940 583520 262340
rect 480 252412 583520 261940
rect 480 252012 583440 252412
rect 480 247380 583520 252012
rect 560 246980 583520 247380
rect 480 240716 583520 246980
rect 480 240316 583440 240716
rect 480 232284 583520 240316
rect 560 231884 583520 232284
rect 480 229020 583520 231884
rect 480 228620 583440 229020
rect 480 217324 583520 228620
rect 560 217188 583520 217324
rect 560 216924 583440 217188
rect 480 216788 583440 216924
rect 480 205492 583520 216788
rect 480 205092 583440 205492
rect 480 202364 583520 205092
rect 560 201964 583520 202364
rect 480 193796 583520 201964
rect 480 193396 583440 193796
rect 480 187404 583520 193396
rect 560 187004 583520 187404
rect 480 182100 583520 187004
rect 480 181700 583440 182100
rect 480 172444 583520 181700
rect 560 172044 583520 172444
rect 480 170268 583520 172044
rect 480 169868 583440 170268
rect 480 158572 583520 169868
rect 480 158172 583440 158572
rect 480 157484 583520 158172
rect 560 157084 583520 157484
rect 480 146876 583520 157084
rect 480 146476 583440 146876
rect 480 142524 583520 146476
rect 560 142124 583520 142524
rect 480 135044 583520 142124
rect 480 134644 583440 135044
rect 480 127564 583520 134644
rect 560 127164 583520 127564
rect 480 123348 583520 127164
rect 480 122948 583440 123348
rect 480 112468 583520 122948
rect 560 112068 583520 112468
rect 480 111652 583520 112068
rect 480 111252 583440 111652
rect 480 99956 583520 111252
rect 480 99556 583440 99956
rect 480 97508 583520 99556
rect 560 97108 583520 97508
rect 480 88124 583520 97108
rect 480 87724 583440 88124
rect 480 82548 583520 87724
rect 560 82148 583520 82548
rect 480 76428 583520 82148
rect 480 76028 583440 76428
rect 480 67588 583520 76028
rect 560 67188 583520 67588
rect 480 64732 583520 67188
rect 480 64332 583440 64732
rect 480 53036 583520 64332
rect 480 52636 583440 53036
rect 480 52628 583520 52636
rect 560 52228 583520 52628
rect 480 41204 583520 52228
rect 480 40804 583440 41204
rect 480 37668 583520 40804
rect 560 37268 583520 37668
rect 480 29508 583520 37268
rect 480 29108 583440 29508
rect 480 22708 583520 29108
rect 560 22308 583520 22708
rect 480 17812 583520 22308
rect 480 17412 583440 17812
rect 480 7748 583520 17412
rect 560 7348 583520 7748
rect 480 6116 583520 7348
rect 480 5716 583440 6116
rect 480 2143 583520 5716
<< metal4 >>
rect -8576 -7504 -7976 711440
rect -7636 -6564 -7036 710500
rect -6696 -5624 -6096 709560
rect -5756 -4684 -5156 708620
rect -4816 -3744 -4216 707680
rect -3876 -2804 -3276 706740
rect -2936 -1864 -2336 705800
rect -1996 -924 -1396 704860
rect 1804 -1864 2404 705800
rect 5404 -3744 6004 707680
rect 9004 -5624 9604 709560
rect 12604 -7504 13204 711440
rect 19804 -1864 20404 705800
rect 23404 -3744 24004 707680
rect 27004 -5624 27604 709560
rect 30604 -7504 31204 711440
rect 37804 -1864 38404 705800
rect 41404 -3744 42004 707680
rect 45004 -5624 45604 709560
rect 48604 -7504 49204 711440
rect 55804 -1864 56404 705800
rect 59404 -3744 60004 707680
rect 63004 -5624 63604 709560
rect 66604 613200 67204 711440
rect 73804 613152 74404 705800
rect 77404 613200 78004 707680
rect 81004 613200 81604 709560
rect 84604 613200 85204 711440
rect 91804 613152 92404 705800
rect 95404 613200 96004 707680
rect 99004 613200 99604 709560
rect 102604 613200 103204 711440
rect 109804 613152 110404 705800
rect 113404 613200 114004 707680
rect 117004 613200 117604 709560
rect 120604 613200 121204 711440
rect 127804 613152 128404 705800
rect 66604 460400 67204 549200
rect 73804 460352 74404 549248
rect 77404 460400 78004 549200
rect 81004 460400 81604 549200
rect 84604 460400 85204 549200
rect 91804 460352 92404 549248
rect 95404 460400 96004 549200
rect 99004 460400 99604 549200
rect 102604 460400 103204 549200
rect 109804 460352 110404 549248
rect 113404 460400 114004 549200
rect 117004 460400 117604 549200
rect 120604 460400 121204 549200
rect 127804 460352 128404 549248
rect 66604 307600 67204 396400
rect 73804 307552 74404 396448
rect 77404 307600 78004 396400
rect 81004 307600 81604 396400
rect 84604 307600 85204 396400
rect 91804 307552 92404 396448
rect 95404 307600 96004 396400
rect 99004 307600 99604 396400
rect 102604 307600 103204 396400
rect 109804 307552 110404 396448
rect 113404 307600 114004 396400
rect 117004 307600 117604 396400
rect 120604 307600 121204 396400
rect 127804 307552 128404 396448
rect 66604 154800 67204 243600
rect 73804 154752 74404 243648
rect 77404 154800 78004 243600
rect 81004 154800 81604 243600
rect 84604 154800 85204 243600
rect 91804 154752 92404 243648
rect 95404 154800 96004 243600
rect 99004 154800 99604 243600
rect 102604 154800 103204 243600
rect 109804 154752 110404 243648
rect 113404 154800 114004 243600
rect 117004 154800 117604 243600
rect 120604 154800 121204 243600
rect 127804 154752 128404 243648
rect 66604 -7504 67204 90800
rect 73804 -1864 74404 90848
rect 77404 -3744 78004 90800
rect 81004 -5624 81604 90800
rect 84604 -7504 85204 90800
rect 91804 -1864 92404 90848
rect 95404 -3744 96004 90800
rect 99004 -5624 99604 90800
rect 102604 -7504 103204 90800
rect 109804 -1864 110404 90848
rect 113404 -3744 114004 90800
rect 117004 -5624 117604 90800
rect 120604 -7504 121204 90800
rect 127804 -1864 128404 90848
rect 131404 -3744 132004 707680
rect 135004 -5624 135604 709560
rect 138604 -7504 139204 711440
rect 145804 -1864 146404 705800
rect 149404 -3744 150004 707680
rect 153004 -5624 153604 709560
rect 156604 -7504 157204 711440
rect 163804 -1864 164404 705800
rect 167404 -3744 168004 707680
rect 171004 -5624 171604 709560
rect 174604 -7504 175204 711440
rect 181804 -1864 182404 705800
rect 185404 -3744 186004 707680
rect 189004 -5624 189604 709560
rect 192604 -7504 193204 711440
rect 199804 613152 200404 705800
rect 203404 613200 204004 707680
rect 207004 613200 207604 709560
rect 210604 613200 211204 711440
rect 217804 613152 218404 705800
rect 221404 613200 222004 707680
rect 225004 613200 225604 709560
rect 228604 613200 229204 711440
rect 235804 613152 236404 705800
rect 239404 613200 240004 707680
rect 243004 613200 243604 709560
rect 246604 613200 247204 711440
rect 253804 613152 254404 705800
rect 257404 613200 258004 707680
rect 199804 460352 200404 549248
rect 203404 460400 204004 549200
rect 207004 460400 207604 549200
rect 210604 460400 211204 549200
rect 217804 460352 218404 549248
rect 221404 460400 222004 549200
rect 225004 460400 225604 549200
rect 228604 460400 229204 549200
rect 235804 460352 236404 549248
rect 239404 460400 240004 549200
rect 243004 460400 243604 549200
rect 246604 460400 247204 549200
rect 253804 460352 254404 549248
rect 257404 460400 258004 549200
rect 199804 307552 200404 396448
rect 203404 307600 204004 396400
rect 207004 307600 207604 396400
rect 210604 307600 211204 396400
rect 217804 307552 218404 396448
rect 221404 307600 222004 396400
rect 225004 307600 225604 396400
rect 228604 307600 229204 396400
rect 235804 307552 236404 396448
rect 239404 307600 240004 396400
rect 243004 307600 243604 396400
rect 246604 307600 247204 396400
rect 253804 307552 254404 396448
rect 257404 307600 258004 396400
rect 199804 154752 200404 243648
rect 203404 154800 204004 243600
rect 207004 154800 207604 243600
rect 210604 154800 211204 243600
rect 217804 154752 218404 243648
rect 221404 154800 222004 243600
rect 225004 154800 225604 243600
rect 228604 154800 229204 243600
rect 235804 154752 236404 243648
rect 239404 154800 240004 243600
rect 243004 154800 243604 243600
rect 246604 154800 247204 243600
rect 253804 154752 254404 243648
rect 257404 154800 258004 243600
rect 199804 -1864 200404 90848
rect 203404 -3744 204004 90800
rect 207004 -5624 207604 90800
rect 210604 -7504 211204 90800
rect 217804 -1864 218404 90848
rect 221404 -3744 222004 90800
rect 225004 -5624 225604 90800
rect 228604 -7504 229204 90800
rect 235804 -1864 236404 90848
rect 239404 -3744 240004 90800
rect 243004 -5624 243604 90800
rect 246604 -7504 247204 90800
rect 253804 -1864 254404 90848
rect 257404 -3744 258004 90800
rect 261004 -5624 261604 709560
rect 264604 -7504 265204 711440
rect 271804 -1864 272404 705800
rect 275404 -3744 276004 707680
rect 279004 -5624 279604 709560
rect 282604 -7504 283204 711440
rect 289804 -1864 290404 705800
rect 293404 -3744 294004 707680
rect 297004 -5624 297604 709560
rect 300604 -7504 301204 711440
rect 307804 -1864 308404 705800
rect 311404 -3744 312004 707680
rect 315004 -5624 315604 709560
rect 318604 -7504 319204 711440
rect 325804 613152 326404 705800
rect 329404 613200 330004 707680
rect 333004 613200 333604 709560
rect 336604 613200 337204 711440
rect 343804 613152 344404 705800
rect 347404 613200 348004 707680
rect 351004 613200 351604 709560
rect 354604 613200 355204 711440
rect 361804 613152 362404 705800
rect 365404 613200 366004 707680
rect 369004 613200 369604 709560
rect 372604 613200 373204 711440
rect 379804 613152 380404 705800
rect 383404 613200 384004 707680
rect 387004 613200 387604 709560
rect 325804 460352 326404 549248
rect 329404 460400 330004 549200
rect 333004 460400 333604 549200
rect 336604 460400 337204 549200
rect 343804 460352 344404 549248
rect 347404 460400 348004 549200
rect 351004 460400 351604 549200
rect 354604 460400 355204 549200
rect 361804 460352 362404 549248
rect 365404 460400 366004 549200
rect 369004 460400 369604 549200
rect 372604 460400 373204 549200
rect 379804 460352 380404 549248
rect 383404 460400 384004 549200
rect 387004 460400 387604 549200
rect 325804 307552 326404 396448
rect 329404 307600 330004 396400
rect 333004 307600 333604 396400
rect 336604 307600 337204 396400
rect 343804 307552 344404 396448
rect 347404 307600 348004 396400
rect 351004 307600 351604 396400
rect 354604 307600 355204 396400
rect 361804 307552 362404 396448
rect 365404 307600 366004 396400
rect 369004 307600 369604 396400
rect 372604 307600 373204 396400
rect 379804 307552 380404 396448
rect 383404 307600 384004 396400
rect 387004 307600 387604 396400
rect 325804 154752 326404 243648
rect 329404 154800 330004 243600
rect 333004 154800 333604 243600
rect 336604 154800 337204 243600
rect 343804 154752 344404 243648
rect 347404 154800 348004 243600
rect 351004 154800 351604 243600
rect 354604 154800 355204 243600
rect 361804 154752 362404 243648
rect 365404 154800 366004 243600
rect 369004 154800 369604 243600
rect 372604 154800 373204 243600
rect 379804 154752 380404 243648
rect 383404 154800 384004 243600
rect 387004 154800 387604 243600
rect 325804 -1864 326404 90848
rect 329404 -3744 330004 90800
rect 333004 -5624 333604 90800
rect 336604 -7504 337204 90800
rect 343804 -1864 344404 90848
rect 347404 -3744 348004 90800
rect 351004 -5624 351604 90800
rect 354604 -7504 355204 90800
rect 361804 -1864 362404 90848
rect 365404 -3744 366004 90800
rect 369004 -5624 369604 90800
rect 372604 -7504 373204 90800
rect 379804 -1864 380404 90848
rect 383404 -3744 384004 90800
rect 387004 -5624 387604 90800
rect 390604 -7504 391204 711440
rect 397804 -1864 398404 705800
rect 401404 -3744 402004 707680
rect 405004 -5624 405604 709560
rect 408604 -7504 409204 711440
rect 415804 -1864 416404 705800
rect 419404 -3744 420004 707680
rect 423004 -5624 423604 709560
rect 426604 -7504 427204 711440
rect 433804 -1864 434404 705800
rect 437404 -3744 438004 707680
rect 441004 -5624 441604 709560
rect 444604 -7504 445204 711440
rect 451804 -1864 452404 705800
rect 455404 613200 456004 707680
rect 459004 613200 459604 709560
rect 462604 613200 463204 711440
rect 469804 613152 470404 705800
rect 473404 613200 474004 707680
rect 477004 613200 477604 709560
rect 480604 613200 481204 711440
rect 487804 613152 488404 705800
rect 491404 613200 492004 707680
rect 495004 613200 495604 709560
rect 498604 613200 499204 711440
rect 505804 613152 506404 705800
rect 509404 613200 510004 707680
rect 513004 613200 513604 709560
rect 516604 613200 517204 711440
rect 455404 460400 456004 549200
rect 459004 460400 459604 549200
rect 462604 460400 463204 549200
rect 469804 460352 470404 549248
rect 473404 460400 474004 549200
rect 477004 460400 477604 549200
rect 480604 460400 481204 549200
rect 487804 460352 488404 549248
rect 491404 460400 492004 549200
rect 495004 460400 495604 549200
rect 498604 460400 499204 549200
rect 505804 460352 506404 549248
rect 509404 460400 510004 549200
rect 513004 460400 513604 549200
rect 516604 460400 517204 549200
rect 455404 307600 456004 396400
rect 459004 307600 459604 396400
rect 462604 307600 463204 396400
rect 469804 307552 470404 396448
rect 473404 307600 474004 396400
rect 477004 307600 477604 396400
rect 480604 307600 481204 396400
rect 487804 307552 488404 396448
rect 491404 307600 492004 396400
rect 495004 307600 495604 396400
rect 498604 307600 499204 396400
rect 505804 307552 506404 396448
rect 509404 307600 510004 396400
rect 513004 307600 513604 396400
rect 516604 307600 517204 396400
rect 455404 154800 456004 243600
rect 459004 154800 459604 243600
rect 462604 154800 463204 243600
rect 469804 154752 470404 243648
rect 473404 154800 474004 243600
rect 477004 154800 477604 243600
rect 480604 154800 481204 243600
rect 487804 154752 488404 243648
rect 491404 154800 492004 243600
rect 495004 154800 495604 243600
rect 498604 154800 499204 243600
rect 505804 154752 506404 243648
rect 509404 154800 510004 243600
rect 513004 154800 513604 243600
rect 516604 154800 517204 243600
rect 455404 -3744 456004 90800
rect 459004 -5624 459604 90800
rect 462604 -7504 463204 90800
rect 469804 -1864 470404 90848
rect 473404 -3744 474004 90800
rect 477004 -5624 477604 90800
rect 480604 -7504 481204 90800
rect 487804 -1864 488404 90848
rect 491404 -3744 492004 90800
rect 495004 -5624 495604 90800
rect 498604 -7504 499204 90800
rect 505804 -1864 506404 90848
rect 509404 -3744 510004 90800
rect 513004 -5624 513604 90800
rect 516604 -7504 517204 90800
rect 523804 -1864 524404 705800
rect 527404 -3744 528004 707680
rect 531004 -5624 531604 709560
rect 534604 -7504 535204 711440
rect 541804 -1864 542404 705800
rect 545404 -3744 546004 707680
rect 549004 -5624 549604 709560
rect 552604 -7504 553204 711440
rect 559804 -1864 560404 705800
rect 563404 -3744 564004 707680
rect 567004 -5624 567604 709560
rect 570604 -7504 571204 711440
rect 577804 -1864 578404 705800
rect 581404 -3744 582004 707680
rect 585320 -924 585920 704860
rect 586260 -1864 586860 705800
rect 587200 -2804 587800 706740
rect 588140 -3744 588740 707680
rect 589080 -4684 589680 708620
rect 590020 -5624 590620 709560
rect 590960 -6564 591560 710500
rect 591900 -7504 592500 711440
<< obsm4 >>
rect 64091 613120 66524 702541
rect 67284 613120 73724 702541
rect 64091 613072 73724 613120
rect 74484 613120 77324 702541
rect 78084 613120 80924 702541
rect 81684 613120 84524 702541
rect 85284 613120 91724 702541
rect 74484 613072 91724 613120
rect 92484 613120 95324 702541
rect 96084 613120 98924 702541
rect 99684 613120 102524 702541
rect 103284 613120 109724 702541
rect 92484 613072 109724 613120
rect 110484 613120 113324 702541
rect 114084 613120 116924 702541
rect 117684 613120 120524 702541
rect 121284 613120 127724 702541
rect 110484 613072 127724 613120
rect 128484 613072 131324 702541
rect 64091 549328 131324 613072
rect 64091 549280 73724 549328
rect 64091 460320 66524 549280
rect 67284 460320 73724 549280
rect 74484 549280 91724 549328
rect 64091 460272 73724 460320
rect 74484 460320 77324 549280
rect 78084 460320 80924 549280
rect 81684 460320 84524 549280
rect 85284 460320 91724 549280
rect 92484 549280 109724 549328
rect 74484 460272 91724 460320
rect 92484 460320 95324 549280
rect 96084 460320 98924 549280
rect 99684 460320 102524 549280
rect 103284 460320 109724 549280
rect 110484 549280 127724 549328
rect 92484 460272 109724 460320
rect 110484 460320 113324 549280
rect 114084 460320 116924 549280
rect 117684 460320 120524 549280
rect 121284 460320 127724 549280
rect 110484 460272 127724 460320
rect 128484 460272 131324 549328
rect 64091 396528 131324 460272
rect 64091 396480 73724 396528
rect 64091 307520 66524 396480
rect 67284 307520 73724 396480
rect 74484 396480 91724 396528
rect 64091 307472 73724 307520
rect 74484 307520 77324 396480
rect 78084 307520 80924 396480
rect 81684 307520 84524 396480
rect 85284 307520 91724 396480
rect 92484 396480 109724 396528
rect 74484 307472 91724 307520
rect 92484 307520 95324 396480
rect 96084 307520 98924 396480
rect 99684 307520 102524 396480
rect 103284 307520 109724 396480
rect 110484 396480 127724 396528
rect 92484 307472 109724 307520
rect 110484 307520 113324 396480
rect 114084 307520 116924 396480
rect 117684 307520 120524 396480
rect 121284 307520 127724 396480
rect 110484 307472 127724 307520
rect 128484 307472 131324 396528
rect 64091 243728 131324 307472
rect 64091 243680 73724 243728
rect 64091 154720 66524 243680
rect 67284 154720 73724 243680
rect 74484 243680 91724 243728
rect 64091 154672 73724 154720
rect 74484 154720 77324 243680
rect 78084 154720 80924 243680
rect 81684 154720 84524 243680
rect 85284 154720 91724 243680
rect 92484 243680 109724 243728
rect 74484 154672 91724 154720
rect 92484 154720 95324 243680
rect 96084 154720 98924 243680
rect 99684 154720 102524 243680
rect 103284 154720 109724 243680
rect 110484 243680 127724 243728
rect 92484 154672 109724 154720
rect 110484 154720 113324 243680
rect 114084 154720 116924 243680
rect 117684 154720 120524 243680
rect 121284 154720 127724 243680
rect 110484 154672 127724 154720
rect 128484 154672 131324 243728
rect 64091 90928 131324 154672
rect 64091 90880 73724 90928
rect 64091 3299 66524 90880
rect 67284 3299 73724 90880
rect 74484 90880 91724 90928
rect 74484 3299 77324 90880
rect 78084 3299 80924 90880
rect 81684 3299 84524 90880
rect 85284 3299 91724 90880
rect 92484 90880 109724 90928
rect 92484 3299 95324 90880
rect 96084 3299 98924 90880
rect 99684 3299 102524 90880
rect 103284 3299 109724 90880
rect 110484 90880 127724 90928
rect 110484 3299 113324 90880
rect 114084 3299 116924 90880
rect 117684 3299 120524 90880
rect 121284 3299 127724 90880
rect 128484 3299 131324 90928
rect 132084 3299 134924 702541
rect 135684 3299 138524 702541
rect 139284 3299 145724 702541
rect 146484 3299 149324 702541
rect 150084 3299 152924 702541
rect 153684 3299 156524 702541
rect 157284 3299 163724 702541
rect 164484 3299 167324 702541
rect 168084 3299 170924 702541
rect 171684 3299 174524 702541
rect 175284 3299 181724 702541
rect 182484 3299 185324 702541
rect 186084 3299 188924 702541
rect 189684 3299 192524 702541
rect 193284 613072 199724 702541
rect 200484 613120 203324 702541
rect 204084 613120 206924 702541
rect 207684 613120 210524 702541
rect 211284 613120 217724 702541
rect 200484 613072 217724 613120
rect 218484 613120 221324 702541
rect 222084 613120 224924 702541
rect 225684 613120 228524 702541
rect 229284 613120 235724 702541
rect 218484 613072 235724 613120
rect 236484 613120 239324 702541
rect 240084 613120 242924 702541
rect 243684 613120 246524 702541
rect 247284 613120 253724 702541
rect 236484 613072 253724 613120
rect 254484 613120 257324 702541
rect 258084 613120 260924 702541
rect 254484 613072 260924 613120
rect 193284 549328 260924 613072
rect 193284 460272 199724 549328
rect 200484 549280 217724 549328
rect 200484 460320 203324 549280
rect 204084 460320 206924 549280
rect 207684 460320 210524 549280
rect 211284 460320 217724 549280
rect 218484 549280 235724 549328
rect 200484 460272 217724 460320
rect 218484 460320 221324 549280
rect 222084 460320 224924 549280
rect 225684 460320 228524 549280
rect 229284 460320 235724 549280
rect 236484 549280 253724 549328
rect 218484 460272 235724 460320
rect 236484 460320 239324 549280
rect 240084 460320 242924 549280
rect 243684 460320 246524 549280
rect 247284 460320 253724 549280
rect 254484 549280 260924 549328
rect 236484 460272 253724 460320
rect 254484 460320 257324 549280
rect 258084 460320 260924 549280
rect 254484 460272 260924 460320
rect 193284 396528 260924 460272
rect 193284 307472 199724 396528
rect 200484 396480 217724 396528
rect 200484 307520 203324 396480
rect 204084 307520 206924 396480
rect 207684 307520 210524 396480
rect 211284 307520 217724 396480
rect 218484 396480 235724 396528
rect 200484 307472 217724 307520
rect 218484 307520 221324 396480
rect 222084 307520 224924 396480
rect 225684 307520 228524 396480
rect 229284 307520 235724 396480
rect 236484 396480 253724 396528
rect 218484 307472 235724 307520
rect 236484 307520 239324 396480
rect 240084 307520 242924 396480
rect 243684 307520 246524 396480
rect 247284 307520 253724 396480
rect 254484 396480 260924 396528
rect 236484 307472 253724 307520
rect 254484 307520 257324 396480
rect 258084 307520 260924 396480
rect 254484 307472 260924 307520
rect 193284 243728 260924 307472
rect 193284 154672 199724 243728
rect 200484 243680 217724 243728
rect 200484 154720 203324 243680
rect 204084 154720 206924 243680
rect 207684 154720 210524 243680
rect 211284 154720 217724 243680
rect 218484 243680 235724 243728
rect 200484 154672 217724 154720
rect 218484 154720 221324 243680
rect 222084 154720 224924 243680
rect 225684 154720 228524 243680
rect 229284 154720 235724 243680
rect 236484 243680 253724 243728
rect 218484 154672 235724 154720
rect 236484 154720 239324 243680
rect 240084 154720 242924 243680
rect 243684 154720 246524 243680
rect 247284 154720 253724 243680
rect 254484 243680 260924 243728
rect 236484 154672 253724 154720
rect 254484 154720 257324 243680
rect 258084 154720 260924 243680
rect 254484 154672 260924 154720
rect 193284 90928 260924 154672
rect 193284 3299 199724 90928
rect 200484 90880 217724 90928
rect 200484 3299 203324 90880
rect 204084 3299 206924 90880
rect 207684 3299 210524 90880
rect 211284 3299 217724 90880
rect 218484 90880 235724 90928
rect 218484 3299 221324 90880
rect 222084 3299 224924 90880
rect 225684 3299 228524 90880
rect 229284 3299 235724 90880
rect 236484 90880 253724 90928
rect 236484 3299 239324 90880
rect 240084 3299 242924 90880
rect 243684 3299 246524 90880
rect 247284 3299 253724 90880
rect 254484 90880 260924 90928
rect 254484 3299 257324 90880
rect 258084 3299 260924 90880
rect 261684 3299 264524 702541
rect 265284 3299 271724 702541
rect 272484 3299 275324 702541
rect 276084 3299 278924 702541
rect 279684 3299 282524 702541
rect 283284 3299 289724 702541
rect 290484 3299 293324 702541
rect 294084 3299 296924 702541
rect 297684 3299 300524 702541
rect 301284 3299 307724 702541
rect 308484 3299 311324 702541
rect 312084 3299 314924 702541
rect 315684 3299 318524 702541
rect 319284 613072 325724 702541
rect 326484 613120 329324 702541
rect 330084 613120 332924 702541
rect 333684 613120 336524 702541
rect 337284 613120 343724 702541
rect 326484 613072 343724 613120
rect 344484 613120 347324 702541
rect 348084 613120 350924 702541
rect 351684 613120 354524 702541
rect 355284 613120 361724 702541
rect 344484 613072 361724 613120
rect 362484 613120 365324 702541
rect 366084 613120 368924 702541
rect 369684 613120 372524 702541
rect 373284 613120 379724 702541
rect 362484 613072 379724 613120
rect 380484 613120 383324 702541
rect 384084 613120 386924 702541
rect 387684 613120 390524 702541
rect 380484 613072 390524 613120
rect 319284 549328 390524 613072
rect 319284 460272 325724 549328
rect 326484 549280 343724 549328
rect 326484 460320 329324 549280
rect 330084 460320 332924 549280
rect 333684 460320 336524 549280
rect 337284 460320 343724 549280
rect 344484 549280 361724 549328
rect 326484 460272 343724 460320
rect 344484 460320 347324 549280
rect 348084 460320 350924 549280
rect 351684 460320 354524 549280
rect 355284 460320 361724 549280
rect 362484 549280 379724 549328
rect 344484 460272 361724 460320
rect 362484 460320 365324 549280
rect 366084 460320 368924 549280
rect 369684 460320 372524 549280
rect 373284 460320 379724 549280
rect 380484 549280 390524 549328
rect 362484 460272 379724 460320
rect 380484 460320 383324 549280
rect 384084 460320 386924 549280
rect 387684 460320 390524 549280
rect 380484 460272 390524 460320
rect 319284 396528 390524 460272
rect 319284 307472 325724 396528
rect 326484 396480 343724 396528
rect 326484 307520 329324 396480
rect 330084 307520 332924 396480
rect 333684 307520 336524 396480
rect 337284 307520 343724 396480
rect 344484 396480 361724 396528
rect 326484 307472 343724 307520
rect 344484 307520 347324 396480
rect 348084 307520 350924 396480
rect 351684 307520 354524 396480
rect 355284 307520 361724 396480
rect 362484 396480 379724 396528
rect 344484 307472 361724 307520
rect 362484 307520 365324 396480
rect 366084 307520 368924 396480
rect 369684 307520 372524 396480
rect 373284 307520 379724 396480
rect 380484 396480 390524 396528
rect 362484 307472 379724 307520
rect 380484 307520 383324 396480
rect 384084 307520 386924 396480
rect 387684 307520 390524 396480
rect 380484 307472 390524 307520
rect 319284 243728 390524 307472
rect 319284 154672 325724 243728
rect 326484 243680 343724 243728
rect 326484 154720 329324 243680
rect 330084 154720 332924 243680
rect 333684 154720 336524 243680
rect 337284 154720 343724 243680
rect 344484 243680 361724 243728
rect 326484 154672 343724 154720
rect 344484 154720 347324 243680
rect 348084 154720 350924 243680
rect 351684 154720 354524 243680
rect 355284 154720 361724 243680
rect 362484 243680 379724 243728
rect 344484 154672 361724 154720
rect 362484 154720 365324 243680
rect 366084 154720 368924 243680
rect 369684 154720 372524 243680
rect 373284 154720 379724 243680
rect 380484 243680 390524 243728
rect 362484 154672 379724 154720
rect 380484 154720 383324 243680
rect 384084 154720 386924 243680
rect 387684 154720 390524 243680
rect 380484 154672 390524 154720
rect 319284 90928 390524 154672
rect 319284 3299 325724 90928
rect 326484 90880 343724 90928
rect 326484 3299 329324 90880
rect 330084 3299 332924 90880
rect 333684 3299 336524 90880
rect 337284 3299 343724 90880
rect 344484 90880 361724 90928
rect 344484 3299 347324 90880
rect 348084 3299 350924 90880
rect 351684 3299 354524 90880
rect 355284 3299 361724 90880
rect 362484 90880 379724 90928
rect 362484 3299 365324 90880
rect 366084 3299 368924 90880
rect 369684 3299 372524 90880
rect 373284 3299 379724 90880
rect 380484 90880 390524 90928
rect 380484 3299 383324 90880
rect 384084 3299 386924 90880
rect 387684 3299 390524 90880
rect 391284 3299 397724 702541
rect 398484 3299 401324 702541
rect 402084 3299 404924 702541
rect 405684 3299 408524 702541
rect 409284 3299 415724 702541
rect 416484 3299 419324 702541
rect 420084 3299 422924 702541
rect 423684 3299 426524 702541
rect 427284 3299 433724 702541
rect 434484 3299 437324 702541
rect 438084 3299 440924 702541
rect 441684 3299 444524 702541
rect 445284 3299 451724 702541
rect 452484 613120 455324 702541
rect 456084 613120 458924 702541
rect 459684 613120 462524 702541
rect 463284 613120 469724 702541
rect 452484 613072 469724 613120
rect 470484 613120 473324 702541
rect 474084 613120 476924 702541
rect 477684 613120 480524 702541
rect 481284 613120 487724 702541
rect 470484 613072 487724 613120
rect 488484 613120 491324 702541
rect 492084 613120 494924 702541
rect 495684 613120 498524 702541
rect 499284 613120 505724 702541
rect 488484 613072 505724 613120
rect 506484 613120 509324 702541
rect 510084 613120 512924 702541
rect 513684 613120 516524 702541
rect 517284 613120 523724 702541
rect 506484 613072 523724 613120
rect 452484 549328 523724 613072
rect 452484 549280 469724 549328
rect 452484 460320 455324 549280
rect 456084 460320 458924 549280
rect 459684 460320 462524 549280
rect 463284 460320 469724 549280
rect 470484 549280 487724 549328
rect 452484 460272 469724 460320
rect 470484 460320 473324 549280
rect 474084 460320 476924 549280
rect 477684 460320 480524 549280
rect 481284 460320 487724 549280
rect 488484 549280 505724 549328
rect 470484 460272 487724 460320
rect 488484 460320 491324 549280
rect 492084 460320 494924 549280
rect 495684 460320 498524 549280
rect 499284 460320 505724 549280
rect 506484 549280 523724 549328
rect 488484 460272 505724 460320
rect 506484 460320 509324 549280
rect 510084 460320 512924 549280
rect 513684 460320 516524 549280
rect 517284 460320 523724 549280
rect 506484 460272 523724 460320
rect 452484 396528 523724 460272
rect 452484 396480 469724 396528
rect 452484 307520 455324 396480
rect 456084 307520 458924 396480
rect 459684 307520 462524 396480
rect 463284 307520 469724 396480
rect 470484 396480 487724 396528
rect 452484 307472 469724 307520
rect 470484 307520 473324 396480
rect 474084 307520 476924 396480
rect 477684 307520 480524 396480
rect 481284 307520 487724 396480
rect 488484 396480 505724 396528
rect 470484 307472 487724 307520
rect 488484 307520 491324 396480
rect 492084 307520 494924 396480
rect 495684 307520 498524 396480
rect 499284 307520 505724 396480
rect 506484 396480 523724 396528
rect 488484 307472 505724 307520
rect 506484 307520 509324 396480
rect 510084 307520 512924 396480
rect 513684 307520 516524 396480
rect 517284 307520 523724 396480
rect 506484 307472 523724 307520
rect 452484 243728 523724 307472
rect 452484 243680 469724 243728
rect 452484 154720 455324 243680
rect 456084 154720 458924 243680
rect 459684 154720 462524 243680
rect 463284 154720 469724 243680
rect 470484 243680 487724 243728
rect 452484 154672 469724 154720
rect 470484 154720 473324 243680
rect 474084 154720 476924 243680
rect 477684 154720 480524 243680
rect 481284 154720 487724 243680
rect 488484 243680 505724 243728
rect 470484 154672 487724 154720
rect 488484 154720 491324 243680
rect 492084 154720 494924 243680
rect 495684 154720 498524 243680
rect 499284 154720 505724 243680
rect 506484 243680 523724 243728
rect 488484 154672 505724 154720
rect 506484 154720 509324 243680
rect 510084 154720 512924 243680
rect 513684 154720 516524 243680
rect 517284 154720 523724 243680
rect 506484 154672 523724 154720
rect 452484 90928 523724 154672
rect 452484 90880 469724 90928
rect 452484 3299 455324 90880
rect 456084 3299 458924 90880
rect 459684 3299 462524 90880
rect 463284 3299 469724 90880
rect 470484 90880 487724 90928
rect 470484 3299 473324 90880
rect 474084 3299 476924 90880
rect 477684 3299 480524 90880
rect 481284 3299 487724 90880
rect 488484 90880 505724 90928
rect 488484 3299 491324 90880
rect 492084 3299 494924 90880
rect 495684 3299 498524 90880
rect 499284 3299 505724 90880
rect 506484 90880 523724 90928
rect 506484 3299 509324 90880
rect 510084 3299 512924 90880
rect 513684 3299 516524 90880
rect 517284 3299 523724 90880
rect 524484 3299 525813 702541
<< metal5 >>
rect -8576 710840 592500 711440
rect -7636 709900 591560 710500
rect -6696 708960 590620 709560
rect -5756 708020 589680 708620
rect -4816 707080 588740 707680
rect -3876 706140 587800 706740
rect -2936 705200 586860 705800
rect -1996 704260 585920 704860
rect -8576 697676 592500 698276
rect -6696 694076 590620 694676
rect -4816 690476 588740 691076
rect -2936 686828 586860 687428
rect -8576 679676 592500 680276
rect -6696 676076 590620 676676
rect -4816 672476 588740 673076
rect -2936 668828 586860 669428
rect -8576 661676 592500 662276
rect -6696 658076 590620 658676
rect -4816 654476 588740 655076
rect -2936 650828 586860 651428
rect -8576 643676 592500 644276
rect -6696 640076 590620 640676
rect -4816 636476 588740 637076
rect -2936 632828 586860 633428
rect -8576 625676 592500 626276
rect -6696 622076 590620 622676
rect -4816 618476 588740 619076
rect -2936 614828 586860 615428
rect -8576 607676 592500 608276
rect -6696 604076 590620 604676
rect -4816 600476 588740 601076
rect -2936 596828 586860 597428
rect -8576 589676 592500 590276
rect -6696 586076 590620 586676
rect -4816 582476 588740 583076
rect -2936 578828 586860 579428
rect -8576 571676 592500 572276
rect -6696 568076 590620 568676
rect -4816 564476 588740 565076
rect -2936 560828 586860 561428
rect -8576 553676 592500 554276
rect -6696 550076 590620 550676
rect -4816 546476 588740 547076
rect -2936 542828 586860 543428
rect -8576 535676 592500 536276
rect -6696 532076 590620 532676
rect -4816 528476 588740 529076
rect -2936 524828 586860 525428
rect -8576 517676 592500 518276
rect -6696 514076 590620 514676
rect -4816 510476 588740 511076
rect -2936 506828 586860 507428
rect -8576 499676 592500 500276
rect -6696 496076 590620 496676
rect -4816 492476 588740 493076
rect -2936 488828 586860 489428
rect -8576 481676 592500 482276
rect -6696 478076 590620 478676
rect -4816 474476 588740 475076
rect -2936 470828 586860 471428
rect -8576 463676 592500 464276
rect -6696 460076 590620 460676
rect -4816 456476 588740 457076
rect -2936 452828 586860 453428
rect -8576 445676 592500 446276
rect -6696 442076 590620 442676
rect -4816 438476 588740 439076
rect -2936 434828 586860 435428
rect -8576 427676 592500 428276
rect -6696 424076 590620 424676
rect -4816 420476 588740 421076
rect -2936 416828 586860 417428
rect -8576 409676 592500 410276
rect -6696 406076 590620 406676
rect -4816 402476 588740 403076
rect -2936 398828 586860 399428
rect -8576 391676 592500 392276
rect -6696 388076 590620 388676
rect -4816 384476 588740 385076
rect -2936 380828 586860 381428
rect -8576 373676 592500 374276
rect -6696 370076 590620 370676
rect -4816 366476 588740 367076
rect -2936 362828 586860 363428
rect -8576 355676 592500 356276
rect -6696 352076 590620 352676
rect -4816 348476 588740 349076
rect -2936 344828 586860 345428
rect -8576 337676 592500 338276
rect -6696 334076 590620 334676
rect -4816 330476 588740 331076
rect -2936 326828 586860 327428
rect -8576 319676 592500 320276
rect -6696 316076 590620 316676
rect -4816 312476 588740 313076
rect -2936 308828 586860 309428
rect -8576 301676 592500 302276
rect -6696 298076 590620 298676
rect -4816 294476 588740 295076
rect -2936 290828 586860 291428
rect -8576 283676 592500 284276
rect -6696 280076 590620 280676
rect -4816 276476 588740 277076
rect -2936 272828 586860 273428
rect -8576 265676 592500 266276
rect -6696 262076 590620 262676
rect -4816 258476 588740 259076
rect -2936 254828 586860 255428
rect -8576 247676 592500 248276
rect -6696 244076 590620 244676
rect -4816 240476 588740 241076
rect -2936 236828 586860 237428
rect -8576 229676 592500 230276
rect -6696 226076 590620 226676
rect -4816 222476 588740 223076
rect -2936 218828 586860 219428
rect -8576 211676 592500 212276
rect -6696 208076 590620 208676
rect -4816 204476 588740 205076
rect -2936 200828 586860 201428
rect -8576 193676 592500 194276
rect -6696 190076 590620 190676
rect -4816 186476 588740 187076
rect -2936 182828 586860 183428
rect -8576 175676 592500 176276
rect -6696 172076 590620 172676
rect -4816 168476 588740 169076
rect -2936 164828 586860 165428
rect -8576 157676 592500 158276
rect -6696 154076 590620 154676
rect -4816 150476 588740 151076
rect -2936 146828 586860 147428
rect -8576 139676 592500 140276
rect -6696 136076 590620 136676
rect -4816 132476 588740 133076
rect -2936 128828 586860 129428
rect -8576 121676 592500 122276
rect -6696 118076 590620 118676
rect -4816 114476 588740 115076
rect -2936 110828 586860 111428
rect -8576 103676 592500 104276
rect -6696 100076 590620 100676
rect -4816 96476 588740 97076
rect -2936 92828 586860 93428
rect -8576 85676 592500 86276
rect -6696 82076 590620 82676
rect -4816 78476 588740 79076
rect -2936 74828 586860 75428
rect -8576 67676 592500 68276
rect -6696 64076 590620 64676
rect -4816 60476 588740 61076
rect -2936 56828 586860 57428
rect -8576 49676 592500 50276
rect -6696 46076 590620 46676
rect -4816 42476 588740 43076
rect -2936 38828 586860 39428
rect -8576 31676 592500 32276
rect -6696 28076 590620 28676
rect -4816 24476 588740 25076
rect -2936 20828 586860 21428
rect -8576 13676 592500 14276
rect -6696 10076 590620 10676
rect -4816 6476 588740 7076
rect -2936 2828 586860 3428
rect -1996 -924 585920 -324
rect -2936 -1864 586860 -1264
rect -3876 -2804 587800 -2204
rect -4816 -3744 588740 -3144
rect -5756 -4684 589680 -4084
rect -6696 -5624 590620 -5024
rect -7636 -6564 591560 -5964
rect -8576 -7504 592500 -6904
<< obsm5 >>
rect -8576 711440 -7976 711442
rect 30604 711440 31204 711442
rect 66604 711440 67204 711442
rect 102604 711440 103204 711442
rect 138604 711440 139204 711442
rect 174604 711440 175204 711442
rect 210604 711440 211204 711442
rect 246604 711440 247204 711442
rect 282604 711440 283204 711442
rect 318604 711440 319204 711442
rect 354604 711440 355204 711442
rect 390604 711440 391204 711442
rect 426604 711440 427204 711442
rect 462604 711440 463204 711442
rect 498604 711440 499204 711442
rect 534604 711440 535204 711442
rect 570604 711440 571204 711442
rect 591900 711440 592500 711442
rect -8576 710838 -7976 710840
rect 30604 710838 31204 710840
rect 66604 710838 67204 710840
rect 102604 710838 103204 710840
rect 138604 710838 139204 710840
rect 174604 710838 175204 710840
rect 210604 710838 211204 710840
rect 246604 710838 247204 710840
rect 282604 710838 283204 710840
rect 318604 710838 319204 710840
rect 354604 710838 355204 710840
rect 390604 710838 391204 710840
rect 426604 710838 427204 710840
rect 462604 710838 463204 710840
rect 498604 710838 499204 710840
rect 534604 710838 535204 710840
rect 570604 710838 571204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 12604 710500 13204 710502
rect 48604 710500 49204 710502
rect 84604 710500 85204 710502
rect 120604 710500 121204 710502
rect 156604 710500 157204 710502
rect 192604 710500 193204 710502
rect 228604 710500 229204 710502
rect 264604 710500 265204 710502
rect 300604 710500 301204 710502
rect 336604 710500 337204 710502
rect 372604 710500 373204 710502
rect 408604 710500 409204 710502
rect 444604 710500 445204 710502
rect 480604 710500 481204 710502
rect 516604 710500 517204 710502
rect 552604 710500 553204 710502
rect 590960 710500 591560 710502
rect -7636 709898 -7036 709900
rect 12604 709898 13204 709900
rect 48604 709898 49204 709900
rect 84604 709898 85204 709900
rect 120604 709898 121204 709900
rect 156604 709898 157204 709900
rect 192604 709898 193204 709900
rect 228604 709898 229204 709900
rect 264604 709898 265204 709900
rect 300604 709898 301204 709900
rect 336604 709898 337204 709900
rect 372604 709898 373204 709900
rect 408604 709898 409204 709900
rect 444604 709898 445204 709900
rect 480604 709898 481204 709900
rect 516604 709898 517204 709900
rect 552604 709898 553204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 27004 709560 27604 709562
rect 63004 709560 63604 709562
rect 99004 709560 99604 709562
rect 135004 709560 135604 709562
rect 171004 709560 171604 709562
rect 207004 709560 207604 709562
rect 243004 709560 243604 709562
rect 279004 709560 279604 709562
rect 315004 709560 315604 709562
rect 351004 709560 351604 709562
rect 387004 709560 387604 709562
rect 423004 709560 423604 709562
rect 459004 709560 459604 709562
rect 495004 709560 495604 709562
rect 531004 709560 531604 709562
rect 567004 709560 567604 709562
rect 590020 709560 590620 709562
rect -6696 708958 -6096 708960
rect 27004 708958 27604 708960
rect 63004 708958 63604 708960
rect 99004 708958 99604 708960
rect 135004 708958 135604 708960
rect 171004 708958 171604 708960
rect 207004 708958 207604 708960
rect 243004 708958 243604 708960
rect 279004 708958 279604 708960
rect 315004 708958 315604 708960
rect 351004 708958 351604 708960
rect 387004 708958 387604 708960
rect 423004 708958 423604 708960
rect 459004 708958 459604 708960
rect 495004 708958 495604 708960
rect 531004 708958 531604 708960
rect 567004 708958 567604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 9004 708620 9604 708622
rect 45004 708620 45604 708622
rect 81004 708620 81604 708622
rect 117004 708620 117604 708622
rect 153004 708620 153604 708622
rect 189004 708620 189604 708622
rect 225004 708620 225604 708622
rect 261004 708620 261604 708622
rect 297004 708620 297604 708622
rect 333004 708620 333604 708622
rect 369004 708620 369604 708622
rect 405004 708620 405604 708622
rect 441004 708620 441604 708622
rect 477004 708620 477604 708622
rect 513004 708620 513604 708622
rect 549004 708620 549604 708622
rect 589080 708620 589680 708622
rect -5756 708018 -5156 708020
rect 9004 708018 9604 708020
rect 45004 708018 45604 708020
rect 81004 708018 81604 708020
rect 117004 708018 117604 708020
rect 153004 708018 153604 708020
rect 189004 708018 189604 708020
rect 225004 708018 225604 708020
rect 261004 708018 261604 708020
rect 297004 708018 297604 708020
rect 333004 708018 333604 708020
rect 369004 708018 369604 708020
rect 405004 708018 405604 708020
rect 441004 708018 441604 708020
rect 477004 708018 477604 708020
rect 513004 708018 513604 708020
rect 549004 708018 549604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 23404 707680 24004 707682
rect 59404 707680 60004 707682
rect 95404 707680 96004 707682
rect 131404 707680 132004 707682
rect 167404 707680 168004 707682
rect 203404 707680 204004 707682
rect 239404 707680 240004 707682
rect 275404 707680 276004 707682
rect 311404 707680 312004 707682
rect 347404 707680 348004 707682
rect 383404 707680 384004 707682
rect 419404 707680 420004 707682
rect 455404 707680 456004 707682
rect 491404 707680 492004 707682
rect 527404 707680 528004 707682
rect 563404 707680 564004 707682
rect 588140 707680 588740 707682
rect -4816 707078 -4216 707080
rect 23404 707078 24004 707080
rect 59404 707078 60004 707080
rect 95404 707078 96004 707080
rect 131404 707078 132004 707080
rect 167404 707078 168004 707080
rect 203404 707078 204004 707080
rect 239404 707078 240004 707080
rect 275404 707078 276004 707080
rect 311404 707078 312004 707080
rect 347404 707078 348004 707080
rect 383404 707078 384004 707080
rect 419404 707078 420004 707080
rect 455404 707078 456004 707080
rect 491404 707078 492004 707080
rect 527404 707078 528004 707080
rect 563404 707078 564004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 5404 706740 6004 706742
rect 41404 706740 42004 706742
rect 77404 706740 78004 706742
rect 113404 706740 114004 706742
rect 149404 706740 150004 706742
rect 185404 706740 186004 706742
rect 221404 706740 222004 706742
rect 257404 706740 258004 706742
rect 293404 706740 294004 706742
rect 329404 706740 330004 706742
rect 365404 706740 366004 706742
rect 401404 706740 402004 706742
rect 437404 706740 438004 706742
rect 473404 706740 474004 706742
rect 509404 706740 510004 706742
rect 545404 706740 546004 706742
rect 581404 706740 582004 706742
rect 587200 706740 587800 706742
rect -3876 706138 -3276 706140
rect 5404 706138 6004 706140
rect 41404 706138 42004 706140
rect 77404 706138 78004 706140
rect 113404 706138 114004 706140
rect 149404 706138 150004 706140
rect 185404 706138 186004 706140
rect 221404 706138 222004 706140
rect 257404 706138 258004 706140
rect 293404 706138 294004 706140
rect 329404 706138 330004 706140
rect 365404 706138 366004 706140
rect 401404 706138 402004 706140
rect 437404 706138 438004 706140
rect 473404 706138 474004 706140
rect 509404 706138 510004 706140
rect 545404 706138 546004 706140
rect 581404 706138 582004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 19804 705800 20404 705802
rect 55804 705800 56404 705802
rect 91804 705800 92404 705802
rect 127804 705800 128404 705802
rect 163804 705800 164404 705802
rect 199804 705800 200404 705802
rect 235804 705800 236404 705802
rect 271804 705800 272404 705802
rect 307804 705800 308404 705802
rect 343804 705800 344404 705802
rect 379804 705800 380404 705802
rect 415804 705800 416404 705802
rect 451804 705800 452404 705802
rect 487804 705800 488404 705802
rect 523804 705800 524404 705802
rect 559804 705800 560404 705802
rect 586260 705800 586860 705802
rect -2936 705198 -2336 705200
rect 19804 705198 20404 705200
rect 55804 705198 56404 705200
rect 91804 705198 92404 705200
rect 127804 705198 128404 705200
rect 163804 705198 164404 705200
rect 199804 705198 200404 705200
rect 235804 705198 236404 705200
rect 271804 705198 272404 705200
rect 307804 705198 308404 705200
rect 343804 705198 344404 705200
rect 379804 705198 380404 705200
rect 415804 705198 416404 705200
rect 451804 705198 452404 705200
rect 487804 705198 488404 705200
rect 523804 705198 524404 705200
rect 559804 705198 560404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 1804 704860 2404 704862
rect 37804 704860 38404 704862
rect 73804 704860 74404 704862
rect 109804 704860 110404 704862
rect 145804 704860 146404 704862
rect 181804 704860 182404 704862
rect 217804 704860 218404 704862
rect 253804 704860 254404 704862
rect 289804 704860 290404 704862
rect 325804 704860 326404 704862
rect 361804 704860 362404 704862
rect 397804 704860 398404 704862
rect 433804 704860 434404 704862
rect 469804 704860 470404 704862
rect 505804 704860 506404 704862
rect 541804 704860 542404 704862
rect 577804 704860 578404 704862
rect 585320 704860 585920 704862
rect -1996 704258 -1396 704260
rect 1804 704258 2404 704260
rect 37804 704258 38404 704260
rect 73804 704258 74404 704260
rect 109804 704258 110404 704260
rect 145804 704258 146404 704260
rect 181804 704258 182404 704260
rect 217804 704258 218404 704260
rect 253804 704258 254404 704260
rect 289804 704258 290404 704260
rect 325804 704258 326404 704260
rect 361804 704258 362404 704260
rect 397804 704258 398404 704260
rect 433804 704258 434404 704260
rect 469804 704258 470404 704260
rect 505804 704258 506404 704260
rect 541804 704258 542404 704260
rect 577804 704258 578404 704260
rect 585320 704258 585920 704260
rect 0 698596 584000 703940
rect -7636 698276 -7036 698278
rect 590960 698276 591560 698278
rect -7636 697674 -7036 697676
rect 590960 697674 591560 697676
rect 0 694996 584000 697356
rect -5756 694676 -5156 694678
rect 589080 694676 589680 694678
rect -5756 694074 -5156 694076
rect 589080 694074 589680 694076
rect 0 691396 584000 693756
rect -3876 691076 -3276 691078
rect 587200 691076 587800 691078
rect -3876 690474 -3276 690476
rect 587200 690474 587800 690476
rect 0 687748 584000 690156
rect -1996 687428 -1396 687430
rect 585320 687428 585920 687430
rect -1996 686826 -1396 686828
rect 585320 686826 585920 686828
rect 0 680596 584000 686508
rect -8576 680276 -7976 680278
rect 591900 680276 592500 680278
rect -8576 679674 -7976 679676
rect 591900 679674 592500 679676
rect 0 676996 584000 679356
rect -6696 676676 -6096 676678
rect 590020 676676 590620 676678
rect -6696 676074 -6096 676076
rect 590020 676074 590620 676076
rect 0 673396 584000 675756
rect -4816 673076 -4216 673078
rect 588140 673076 588740 673078
rect -4816 672474 -4216 672476
rect 588140 672474 588740 672476
rect 0 669748 584000 672156
rect -2936 669428 -2336 669430
rect 586260 669428 586860 669430
rect -2936 668826 -2336 668828
rect 586260 668826 586860 668828
rect 0 662596 584000 668508
rect -7636 662276 -7036 662278
rect 590960 662276 591560 662278
rect -7636 661674 -7036 661676
rect 590960 661674 591560 661676
rect 0 658996 584000 661356
rect -5756 658676 -5156 658678
rect 589080 658676 589680 658678
rect -5756 658074 -5156 658076
rect 589080 658074 589680 658076
rect 0 655396 584000 657756
rect -3876 655076 -3276 655078
rect 587200 655076 587800 655078
rect -3876 654474 -3276 654476
rect 587200 654474 587800 654476
rect 0 651748 584000 654156
rect -1996 651428 -1396 651430
rect 585320 651428 585920 651430
rect -1996 650826 -1396 650828
rect 585320 650826 585920 650828
rect 0 644596 584000 650508
rect -8576 644276 -7976 644278
rect 591900 644276 592500 644278
rect -8576 643674 -7976 643676
rect 591900 643674 592500 643676
rect 0 640996 584000 643356
rect -6696 640676 -6096 640678
rect 590020 640676 590620 640678
rect -6696 640074 -6096 640076
rect 590020 640074 590620 640076
rect 0 637396 584000 639756
rect -4816 637076 -4216 637078
rect 588140 637076 588740 637078
rect -4816 636474 -4216 636476
rect 588140 636474 588740 636476
rect 0 633748 584000 636156
rect -2936 633428 -2336 633430
rect 586260 633428 586860 633430
rect -2936 632826 -2336 632828
rect 586260 632826 586860 632828
rect 0 626596 584000 632508
rect -7636 626276 -7036 626278
rect 590960 626276 591560 626278
rect -7636 625674 -7036 625676
rect 590960 625674 591560 625676
rect 0 622996 584000 625356
rect -5756 622676 -5156 622678
rect 589080 622676 589680 622678
rect -5756 622074 -5156 622076
rect 589080 622074 589680 622076
rect 0 619396 584000 621756
rect -3876 619076 -3276 619078
rect 587200 619076 587800 619078
rect -3876 618474 -3276 618476
rect 587200 618474 587800 618476
rect 0 615748 584000 618156
rect -1996 615428 -1396 615430
rect 585320 615428 585920 615430
rect -1996 614826 -1396 614828
rect 585320 614826 585920 614828
rect 0 608596 584000 614508
rect -8576 608276 -7976 608278
rect 591900 608276 592500 608278
rect -8576 607674 -7976 607676
rect 591900 607674 592500 607676
rect 0 604996 584000 607356
rect -6696 604676 -6096 604678
rect 590020 604676 590620 604678
rect -6696 604074 -6096 604076
rect 590020 604074 590620 604076
rect 0 601396 584000 603756
rect -4816 601076 -4216 601078
rect 588140 601076 588740 601078
rect -4816 600474 -4216 600476
rect 588140 600474 588740 600476
rect 0 597748 584000 600156
rect -2936 597428 -2336 597430
rect 586260 597428 586860 597430
rect -2936 596826 -2336 596828
rect 586260 596826 586860 596828
rect 0 590596 584000 596508
rect -7636 590276 -7036 590278
rect 590960 590276 591560 590278
rect -7636 589674 -7036 589676
rect 590960 589674 591560 589676
rect 0 586996 584000 589356
rect -5756 586676 -5156 586678
rect 589080 586676 589680 586678
rect -5756 586074 -5156 586076
rect 589080 586074 589680 586076
rect 0 583396 584000 585756
rect -3876 583076 -3276 583078
rect 587200 583076 587800 583078
rect -3876 582474 -3276 582476
rect 587200 582474 587800 582476
rect 0 579748 584000 582156
rect -1996 579428 -1396 579430
rect 585320 579428 585920 579430
rect -1996 578826 -1396 578828
rect 585320 578826 585920 578828
rect 0 572596 584000 578508
rect -8576 572276 -7976 572278
rect 591900 572276 592500 572278
rect -8576 571674 -7976 571676
rect 591900 571674 592500 571676
rect 0 568996 584000 571356
rect -6696 568676 -6096 568678
rect 590020 568676 590620 568678
rect -6696 568074 -6096 568076
rect 590020 568074 590620 568076
rect 0 565396 584000 567756
rect -4816 565076 -4216 565078
rect 588140 565076 588740 565078
rect -4816 564474 -4216 564476
rect 588140 564474 588740 564476
rect 0 561748 584000 564156
rect -2936 561428 -2336 561430
rect 586260 561428 586860 561430
rect -2936 560826 -2336 560828
rect 586260 560826 586860 560828
rect 0 554596 584000 560508
rect -7636 554276 -7036 554278
rect 590960 554276 591560 554278
rect -7636 553674 -7036 553676
rect 590960 553674 591560 553676
rect 0 550996 584000 553356
rect -5756 550676 -5156 550678
rect 589080 550676 589680 550678
rect -5756 550074 -5156 550076
rect 589080 550074 589680 550076
rect 0 547396 584000 549756
rect -3876 547076 -3276 547078
rect 587200 547076 587800 547078
rect -3876 546474 -3276 546476
rect 587200 546474 587800 546476
rect 0 543748 584000 546156
rect -1996 543428 -1396 543430
rect 585320 543428 585920 543430
rect -1996 542826 -1396 542828
rect 585320 542826 585920 542828
rect 0 536596 584000 542508
rect -8576 536276 -7976 536278
rect 591900 536276 592500 536278
rect -8576 535674 -7976 535676
rect 591900 535674 592500 535676
rect 0 532996 584000 535356
rect -6696 532676 -6096 532678
rect 590020 532676 590620 532678
rect -6696 532074 -6096 532076
rect 590020 532074 590620 532076
rect 0 529396 584000 531756
rect -4816 529076 -4216 529078
rect 588140 529076 588740 529078
rect -4816 528474 -4216 528476
rect 588140 528474 588740 528476
rect 0 525748 584000 528156
rect -2936 525428 -2336 525430
rect 586260 525428 586860 525430
rect -2936 524826 -2336 524828
rect 586260 524826 586860 524828
rect 0 518596 584000 524508
rect -7636 518276 -7036 518278
rect 590960 518276 591560 518278
rect -7636 517674 -7036 517676
rect 590960 517674 591560 517676
rect 0 514996 584000 517356
rect -5756 514676 -5156 514678
rect 589080 514676 589680 514678
rect -5756 514074 -5156 514076
rect 589080 514074 589680 514076
rect 0 511396 584000 513756
rect -3876 511076 -3276 511078
rect 587200 511076 587800 511078
rect -3876 510474 -3276 510476
rect 587200 510474 587800 510476
rect 0 507748 584000 510156
rect -1996 507428 -1396 507430
rect 585320 507428 585920 507430
rect -1996 506826 -1396 506828
rect 585320 506826 585920 506828
rect 0 500596 584000 506508
rect -8576 500276 -7976 500278
rect 591900 500276 592500 500278
rect -8576 499674 -7976 499676
rect 591900 499674 592500 499676
rect 0 496996 584000 499356
rect -6696 496676 -6096 496678
rect 590020 496676 590620 496678
rect -6696 496074 -6096 496076
rect 590020 496074 590620 496076
rect 0 493396 584000 495756
rect -4816 493076 -4216 493078
rect 588140 493076 588740 493078
rect -4816 492474 -4216 492476
rect 588140 492474 588740 492476
rect 0 489748 584000 492156
rect -2936 489428 -2336 489430
rect 586260 489428 586860 489430
rect -2936 488826 -2336 488828
rect 586260 488826 586860 488828
rect 0 482596 584000 488508
rect -7636 482276 -7036 482278
rect 590960 482276 591560 482278
rect -7636 481674 -7036 481676
rect 590960 481674 591560 481676
rect 0 478996 584000 481356
rect -5756 478676 -5156 478678
rect 589080 478676 589680 478678
rect -5756 478074 -5156 478076
rect 589080 478074 589680 478076
rect 0 475396 584000 477756
rect -3876 475076 -3276 475078
rect 587200 475076 587800 475078
rect -3876 474474 -3276 474476
rect 587200 474474 587800 474476
rect 0 471748 584000 474156
rect -1996 471428 -1396 471430
rect 585320 471428 585920 471430
rect -1996 470826 -1396 470828
rect 585320 470826 585920 470828
rect 0 464596 584000 470508
rect -8576 464276 -7976 464278
rect 591900 464276 592500 464278
rect -8576 463674 -7976 463676
rect 591900 463674 592500 463676
rect 0 460996 584000 463356
rect -6696 460676 -6096 460678
rect 590020 460676 590620 460678
rect -6696 460074 -6096 460076
rect 590020 460074 590620 460076
rect 0 457396 584000 459756
rect -4816 457076 -4216 457078
rect 588140 457076 588740 457078
rect -4816 456474 -4216 456476
rect 588140 456474 588740 456476
rect 0 453748 584000 456156
rect -2936 453428 -2336 453430
rect 586260 453428 586860 453430
rect -2936 452826 -2336 452828
rect 586260 452826 586860 452828
rect 0 446596 584000 452508
rect -7636 446276 -7036 446278
rect 590960 446276 591560 446278
rect -7636 445674 -7036 445676
rect 590960 445674 591560 445676
rect 0 442996 584000 445356
rect -5756 442676 -5156 442678
rect 589080 442676 589680 442678
rect -5756 442074 -5156 442076
rect 589080 442074 589680 442076
rect 0 439396 584000 441756
rect -3876 439076 -3276 439078
rect 587200 439076 587800 439078
rect -3876 438474 -3276 438476
rect 587200 438474 587800 438476
rect 0 435748 584000 438156
rect -1996 435428 -1396 435430
rect 585320 435428 585920 435430
rect -1996 434826 -1396 434828
rect 585320 434826 585920 434828
rect 0 428596 584000 434508
rect -8576 428276 -7976 428278
rect 591900 428276 592500 428278
rect -8576 427674 -7976 427676
rect 591900 427674 592500 427676
rect 0 424996 584000 427356
rect -6696 424676 -6096 424678
rect 590020 424676 590620 424678
rect -6696 424074 -6096 424076
rect 590020 424074 590620 424076
rect 0 421396 584000 423756
rect -4816 421076 -4216 421078
rect 588140 421076 588740 421078
rect -4816 420474 -4216 420476
rect 588140 420474 588740 420476
rect 0 417748 584000 420156
rect -2936 417428 -2336 417430
rect 586260 417428 586860 417430
rect -2936 416826 -2336 416828
rect 586260 416826 586860 416828
rect 0 410596 584000 416508
rect -7636 410276 -7036 410278
rect 590960 410276 591560 410278
rect -7636 409674 -7036 409676
rect 590960 409674 591560 409676
rect 0 406996 584000 409356
rect -5756 406676 -5156 406678
rect 589080 406676 589680 406678
rect -5756 406074 -5156 406076
rect 589080 406074 589680 406076
rect 0 403396 584000 405756
rect -3876 403076 -3276 403078
rect 587200 403076 587800 403078
rect -3876 402474 -3276 402476
rect 587200 402474 587800 402476
rect 0 399748 584000 402156
rect -1996 399428 -1396 399430
rect 585320 399428 585920 399430
rect -1996 398826 -1396 398828
rect 585320 398826 585920 398828
rect 0 392596 584000 398508
rect -8576 392276 -7976 392278
rect 591900 392276 592500 392278
rect -8576 391674 -7976 391676
rect 591900 391674 592500 391676
rect 0 388996 584000 391356
rect -6696 388676 -6096 388678
rect 590020 388676 590620 388678
rect -6696 388074 -6096 388076
rect 590020 388074 590620 388076
rect 0 385396 584000 387756
rect -4816 385076 -4216 385078
rect 588140 385076 588740 385078
rect -4816 384474 -4216 384476
rect 588140 384474 588740 384476
rect 0 381748 584000 384156
rect -2936 381428 -2336 381430
rect 586260 381428 586860 381430
rect -2936 380826 -2336 380828
rect 586260 380826 586860 380828
rect 0 374596 584000 380508
rect -7636 374276 -7036 374278
rect 590960 374276 591560 374278
rect -7636 373674 -7036 373676
rect 590960 373674 591560 373676
rect 0 370996 584000 373356
rect -5756 370676 -5156 370678
rect 589080 370676 589680 370678
rect -5756 370074 -5156 370076
rect 589080 370074 589680 370076
rect 0 367396 584000 369756
rect -3876 367076 -3276 367078
rect 587200 367076 587800 367078
rect -3876 366474 -3276 366476
rect 587200 366474 587800 366476
rect 0 363748 584000 366156
rect -1996 363428 -1396 363430
rect 585320 363428 585920 363430
rect -1996 362826 -1396 362828
rect 585320 362826 585920 362828
rect 0 356596 584000 362508
rect -8576 356276 -7976 356278
rect 591900 356276 592500 356278
rect -8576 355674 -7976 355676
rect 591900 355674 592500 355676
rect 0 352996 584000 355356
rect -6696 352676 -6096 352678
rect 590020 352676 590620 352678
rect -6696 352074 -6096 352076
rect 590020 352074 590620 352076
rect 0 349396 584000 351756
rect -4816 349076 -4216 349078
rect 588140 349076 588740 349078
rect -4816 348474 -4216 348476
rect 588140 348474 588740 348476
rect 0 345748 584000 348156
rect -2936 345428 -2336 345430
rect 586260 345428 586860 345430
rect -2936 344826 -2336 344828
rect 586260 344826 586860 344828
rect 0 338596 584000 344508
rect -7636 338276 -7036 338278
rect 590960 338276 591560 338278
rect -7636 337674 -7036 337676
rect 590960 337674 591560 337676
rect 0 334996 584000 337356
rect -5756 334676 -5156 334678
rect 589080 334676 589680 334678
rect -5756 334074 -5156 334076
rect 589080 334074 589680 334076
rect 0 331396 584000 333756
rect -3876 331076 -3276 331078
rect 587200 331076 587800 331078
rect -3876 330474 -3276 330476
rect 587200 330474 587800 330476
rect 0 327748 584000 330156
rect -1996 327428 -1396 327430
rect 585320 327428 585920 327430
rect -1996 326826 -1396 326828
rect 585320 326826 585920 326828
rect 0 320596 584000 326508
rect -8576 320276 -7976 320278
rect 591900 320276 592500 320278
rect -8576 319674 -7976 319676
rect 591900 319674 592500 319676
rect 0 316996 584000 319356
rect -6696 316676 -6096 316678
rect 590020 316676 590620 316678
rect -6696 316074 -6096 316076
rect 590020 316074 590620 316076
rect 0 313396 584000 315756
rect -4816 313076 -4216 313078
rect 588140 313076 588740 313078
rect -4816 312474 -4216 312476
rect 588140 312474 588740 312476
rect 0 309748 584000 312156
rect -2936 309428 -2336 309430
rect 586260 309428 586860 309430
rect -2936 308826 -2336 308828
rect 586260 308826 586860 308828
rect 0 302596 584000 308508
rect -7636 302276 -7036 302278
rect 590960 302276 591560 302278
rect -7636 301674 -7036 301676
rect 590960 301674 591560 301676
rect 0 298996 584000 301356
rect -5756 298676 -5156 298678
rect 589080 298676 589680 298678
rect -5756 298074 -5156 298076
rect 589080 298074 589680 298076
rect 0 295396 584000 297756
rect -3876 295076 -3276 295078
rect 587200 295076 587800 295078
rect -3876 294474 -3276 294476
rect 587200 294474 587800 294476
rect 0 291748 584000 294156
rect -1996 291428 -1396 291430
rect 585320 291428 585920 291430
rect -1996 290826 -1396 290828
rect 585320 290826 585920 290828
rect 0 284596 584000 290508
rect -8576 284276 -7976 284278
rect 591900 284276 592500 284278
rect -8576 283674 -7976 283676
rect 591900 283674 592500 283676
rect 0 280996 584000 283356
rect -6696 280676 -6096 280678
rect 590020 280676 590620 280678
rect -6696 280074 -6096 280076
rect 590020 280074 590620 280076
rect 0 277396 584000 279756
rect -4816 277076 -4216 277078
rect 588140 277076 588740 277078
rect -4816 276474 -4216 276476
rect 588140 276474 588740 276476
rect 0 273748 584000 276156
rect -2936 273428 -2336 273430
rect 586260 273428 586860 273430
rect -2936 272826 -2336 272828
rect 586260 272826 586860 272828
rect 0 266596 584000 272508
rect -7636 266276 -7036 266278
rect 590960 266276 591560 266278
rect -7636 265674 -7036 265676
rect 590960 265674 591560 265676
rect 0 262996 584000 265356
rect -5756 262676 -5156 262678
rect 589080 262676 589680 262678
rect -5756 262074 -5156 262076
rect 589080 262074 589680 262076
rect 0 259396 584000 261756
rect -3876 259076 -3276 259078
rect 587200 259076 587800 259078
rect -3876 258474 -3276 258476
rect 587200 258474 587800 258476
rect 0 255748 584000 258156
rect -1996 255428 -1396 255430
rect 585320 255428 585920 255430
rect -1996 254826 -1396 254828
rect 585320 254826 585920 254828
rect 0 248596 584000 254508
rect -8576 248276 -7976 248278
rect 591900 248276 592500 248278
rect -8576 247674 -7976 247676
rect 591900 247674 592500 247676
rect 0 244996 584000 247356
rect -6696 244676 -6096 244678
rect 590020 244676 590620 244678
rect -6696 244074 -6096 244076
rect 590020 244074 590620 244076
rect 0 241396 584000 243756
rect -4816 241076 -4216 241078
rect 588140 241076 588740 241078
rect -4816 240474 -4216 240476
rect 588140 240474 588740 240476
rect 0 237748 584000 240156
rect -2936 237428 -2336 237430
rect 586260 237428 586860 237430
rect -2936 236826 -2336 236828
rect 586260 236826 586860 236828
rect 0 230596 584000 236508
rect -7636 230276 -7036 230278
rect 590960 230276 591560 230278
rect -7636 229674 -7036 229676
rect 590960 229674 591560 229676
rect 0 226996 584000 229356
rect -5756 226676 -5156 226678
rect 589080 226676 589680 226678
rect -5756 226074 -5156 226076
rect 589080 226074 589680 226076
rect 0 223396 584000 225756
rect -3876 223076 -3276 223078
rect 587200 223076 587800 223078
rect -3876 222474 -3276 222476
rect 587200 222474 587800 222476
rect 0 219748 584000 222156
rect -1996 219428 -1396 219430
rect 585320 219428 585920 219430
rect -1996 218826 -1396 218828
rect 585320 218826 585920 218828
rect 0 212596 584000 218508
rect -8576 212276 -7976 212278
rect 591900 212276 592500 212278
rect -8576 211674 -7976 211676
rect 591900 211674 592500 211676
rect 0 208996 584000 211356
rect -6696 208676 -6096 208678
rect 590020 208676 590620 208678
rect -6696 208074 -6096 208076
rect 590020 208074 590620 208076
rect 0 205396 584000 207756
rect -4816 205076 -4216 205078
rect 588140 205076 588740 205078
rect -4816 204474 -4216 204476
rect 588140 204474 588740 204476
rect 0 201748 584000 204156
rect -2936 201428 -2336 201430
rect 586260 201428 586860 201430
rect -2936 200826 -2336 200828
rect 586260 200826 586860 200828
rect 0 194596 584000 200508
rect -7636 194276 -7036 194278
rect 590960 194276 591560 194278
rect -7636 193674 -7036 193676
rect 590960 193674 591560 193676
rect 0 190996 584000 193356
rect -5756 190676 -5156 190678
rect 589080 190676 589680 190678
rect -5756 190074 -5156 190076
rect 589080 190074 589680 190076
rect 0 187396 584000 189756
rect -3876 187076 -3276 187078
rect 587200 187076 587800 187078
rect -3876 186474 -3276 186476
rect 587200 186474 587800 186476
rect 0 183748 584000 186156
rect -1996 183428 -1396 183430
rect 585320 183428 585920 183430
rect -1996 182826 -1396 182828
rect 585320 182826 585920 182828
rect 0 176596 584000 182508
rect -8576 176276 -7976 176278
rect 591900 176276 592500 176278
rect -8576 175674 -7976 175676
rect 591900 175674 592500 175676
rect 0 172996 584000 175356
rect -6696 172676 -6096 172678
rect 590020 172676 590620 172678
rect -6696 172074 -6096 172076
rect 590020 172074 590620 172076
rect 0 169396 584000 171756
rect -4816 169076 -4216 169078
rect 588140 169076 588740 169078
rect -4816 168474 -4216 168476
rect 588140 168474 588740 168476
rect 0 165748 584000 168156
rect -2936 165428 -2336 165430
rect 586260 165428 586860 165430
rect -2936 164826 -2336 164828
rect 586260 164826 586860 164828
rect 0 158596 584000 164508
rect -7636 158276 -7036 158278
rect 590960 158276 591560 158278
rect -7636 157674 -7036 157676
rect 590960 157674 591560 157676
rect 0 154996 584000 157356
rect -5756 154676 -5156 154678
rect 589080 154676 589680 154678
rect -5756 154074 -5156 154076
rect 589080 154074 589680 154076
rect 0 151396 584000 153756
rect -3876 151076 -3276 151078
rect 587200 151076 587800 151078
rect -3876 150474 -3276 150476
rect 587200 150474 587800 150476
rect 0 147748 584000 150156
rect -1996 147428 -1396 147430
rect 585320 147428 585920 147430
rect -1996 146826 -1396 146828
rect 585320 146826 585920 146828
rect 0 140596 584000 146508
rect -8576 140276 -7976 140278
rect 591900 140276 592500 140278
rect -8576 139674 -7976 139676
rect 591900 139674 592500 139676
rect 0 136996 584000 139356
rect -6696 136676 -6096 136678
rect 590020 136676 590620 136678
rect -6696 136074 -6096 136076
rect 590020 136074 590620 136076
rect 0 133396 584000 135756
rect -4816 133076 -4216 133078
rect 588140 133076 588740 133078
rect -4816 132474 -4216 132476
rect 588140 132474 588740 132476
rect 0 129748 584000 132156
rect -2936 129428 -2336 129430
rect 586260 129428 586860 129430
rect -2936 128826 -2336 128828
rect 586260 128826 586860 128828
rect 0 122596 584000 128508
rect -7636 122276 -7036 122278
rect 590960 122276 591560 122278
rect -7636 121674 -7036 121676
rect 590960 121674 591560 121676
rect 0 118996 584000 121356
rect -5756 118676 -5156 118678
rect 589080 118676 589680 118678
rect -5756 118074 -5156 118076
rect 589080 118074 589680 118076
rect 0 115396 584000 117756
rect -3876 115076 -3276 115078
rect 587200 115076 587800 115078
rect -3876 114474 -3276 114476
rect 587200 114474 587800 114476
rect 0 111748 584000 114156
rect -1996 111428 -1396 111430
rect 585320 111428 585920 111430
rect -1996 110826 -1396 110828
rect 585320 110826 585920 110828
rect 0 104596 584000 110508
rect -8576 104276 -7976 104278
rect 591900 104276 592500 104278
rect -8576 103674 -7976 103676
rect 591900 103674 592500 103676
rect 0 100996 584000 103356
rect -6696 100676 -6096 100678
rect 590020 100676 590620 100678
rect -6696 100074 -6096 100076
rect 590020 100074 590620 100076
rect 0 97396 584000 99756
rect -4816 97076 -4216 97078
rect 588140 97076 588740 97078
rect -4816 96474 -4216 96476
rect 588140 96474 588740 96476
rect 0 93748 584000 96156
rect -2936 93428 -2336 93430
rect 586260 93428 586860 93430
rect -2936 92826 -2336 92828
rect 586260 92826 586860 92828
rect 0 86596 584000 92508
rect -7636 86276 -7036 86278
rect 590960 86276 591560 86278
rect -7636 85674 -7036 85676
rect 590960 85674 591560 85676
rect 0 82996 584000 85356
rect -5756 82676 -5156 82678
rect 589080 82676 589680 82678
rect -5756 82074 -5156 82076
rect 589080 82074 589680 82076
rect 0 79396 584000 81756
rect -3876 79076 -3276 79078
rect 587200 79076 587800 79078
rect -3876 78474 -3276 78476
rect 587200 78474 587800 78476
rect 0 75748 584000 78156
rect -1996 75428 -1396 75430
rect 585320 75428 585920 75430
rect -1996 74826 -1396 74828
rect 585320 74826 585920 74828
rect 0 68596 584000 74508
rect -8576 68276 -7976 68278
rect 591900 68276 592500 68278
rect -8576 67674 -7976 67676
rect 591900 67674 592500 67676
rect 0 64996 584000 67356
rect -6696 64676 -6096 64678
rect 590020 64676 590620 64678
rect -6696 64074 -6096 64076
rect 590020 64074 590620 64076
rect 0 61396 584000 63756
rect -4816 61076 -4216 61078
rect 588140 61076 588740 61078
rect -4816 60474 -4216 60476
rect 588140 60474 588740 60476
rect 0 57748 584000 60156
rect -2936 57428 -2336 57430
rect 586260 57428 586860 57430
rect -2936 56826 -2336 56828
rect 586260 56826 586860 56828
rect 0 50596 584000 56508
rect -7636 50276 -7036 50278
rect 590960 50276 591560 50278
rect -7636 49674 -7036 49676
rect 590960 49674 591560 49676
rect 0 46996 584000 49356
rect -5756 46676 -5156 46678
rect 589080 46676 589680 46678
rect -5756 46074 -5156 46076
rect 589080 46074 589680 46076
rect 0 43396 584000 45756
rect -3876 43076 -3276 43078
rect 587200 43076 587800 43078
rect -3876 42474 -3276 42476
rect 587200 42474 587800 42476
rect 0 39748 584000 42156
rect -1996 39428 -1396 39430
rect 585320 39428 585920 39430
rect -1996 38826 -1396 38828
rect 585320 38826 585920 38828
rect 0 32596 584000 38508
rect -8576 32276 -7976 32278
rect 591900 32276 592500 32278
rect -8576 31674 -7976 31676
rect 591900 31674 592500 31676
rect 0 28996 584000 31356
rect -6696 28676 -6096 28678
rect 590020 28676 590620 28678
rect -6696 28074 -6096 28076
rect 590020 28074 590620 28076
rect 0 25396 584000 27756
rect -4816 25076 -4216 25078
rect 588140 25076 588740 25078
rect -4816 24474 -4216 24476
rect 588140 24474 588740 24476
rect 0 21748 584000 24156
rect -2936 21428 -2336 21430
rect 586260 21428 586860 21430
rect -2936 20826 -2336 20828
rect 586260 20826 586860 20828
rect 0 14596 584000 20508
rect -7636 14276 -7036 14278
rect 590960 14276 591560 14278
rect -7636 13674 -7036 13676
rect 590960 13674 591560 13676
rect 0 10996 584000 13356
rect -5756 10676 -5156 10678
rect 589080 10676 589680 10678
rect -5756 10074 -5156 10076
rect 589080 10074 589680 10076
rect 0 7396 584000 9756
rect -3876 7076 -3276 7078
rect 587200 7076 587800 7078
rect -3876 6474 -3276 6476
rect 587200 6474 587800 6476
rect 0 3748 584000 6156
rect -1996 3428 -1396 3430
rect 585320 3428 585920 3430
rect -1996 2826 -1396 2828
rect 585320 2826 585920 2828
rect 0 0 584000 2508
rect -1996 -324 -1396 -322
rect 1804 -324 2404 -322
rect 37804 -324 38404 -322
rect 73804 -324 74404 -322
rect 109804 -324 110404 -322
rect 145804 -324 146404 -322
rect 181804 -324 182404 -322
rect 217804 -324 218404 -322
rect 253804 -324 254404 -322
rect 289804 -324 290404 -322
rect 325804 -324 326404 -322
rect 361804 -324 362404 -322
rect 397804 -324 398404 -322
rect 433804 -324 434404 -322
rect 469804 -324 470404 -322
rect 505804 -324 506404 -322
rect 541804 -324 542404 -322
rect 577804 -324 578404 -322
rect 585320 -324 585920 -322
rect -1996 -926 -1396 -924
rect 1804 -926 2404 -924
rect 37804 -926 38404 -924
rect 73804 -926 74404 -924
rect 109804 -926 110404 -924
rect 145804 -926 146404 -924
rect 181804 -926 182404 -924
rect 217804 -926 218404 -924
rect 253804 -926 254404 -924
rect 289804 -926 290404 -924
rect 325804 -926 326404 -924
rect 361804 -926 362404 -924
rect 397804 -926 398404 -924
rect 433804 -926 434404 -924
rect 469804 -926 470404 -924
rect 505804 -926 506404 -924
rect 541804 -926 542404 -924
rect 577804 -926 578404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 19804 -1264 20404 -1262
rect 55804 -1264 56404 -1262
rect 91804 -1264 92404 -1262
rect 127804 -1264 128404 -1262
rect 163804 -1264 164404 -1262
rect 199804 -1264 200404 -1262
rect 235804 -1264 236404 -1262
rect 271804 -1264 272404 -1262
rect 307804 -1264 308404 -1262
rect 343804 -1264 344404 -1262
rect 379804 -1264 380404 -1262
rect 415804 -1264 416404 -1262
rect 451804 -1264 452404 -1262
rect 487804 -1264 488404 -1262
rect 523804 -1264 524404 -1262
rect 559804 -1264 560404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1866 -2336 -1864
rect 19804 -1866 20404 -1864
rect 55804 -1866 56404 -1864
rect 91804 -1866 92404 -1864
rect 127804 -1866 128404 -1864
rect 163804 -1866 164404 -1864
rect 199804 -1866 200404 -1864
rect 235804 -1866 236404 -1864
rect 271804 -1866 272404 -1864
rect 307804 -1866 308404 -1864
rect 343804 -1866 344404 -1864
rect 379804 -1866 380404 -1864
rect 415804 -1866 416404 -1864
rect 451804 -1866 452404 -1864
rect 487804 -1866 488404 -1864
rect 523804 -1866 524404 -1864
rect 559804 -1866 560404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 5404 -2204 6004 -2202
rect 41404 -2204 42004 -2202
rect 77404 -2204 78004 -2202
rect 113404 -2204 114004 -2202
rect 149404 -2204 150004 -2202
rect 185404 -2204 186004 -2202
rect 221404 -2204 222004 -2202
rect 257404 -2204 258004 -2202
rect 293404 -2204 294004 -2202
rect 329404 -2204 330004 -2202
rect 365404 -2204 366004 -2202
rect 401404 -2204 402004 -2202
rect 437404 -2204 438004 -2202
rect 473404 -2204 474004 -2202
rect 509404 -2204 510004 -2202
rect 545404 -2204 546004 -2202
rect 581404 -2204 582004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2806 -3276 -2804
rect 5404 -2806 6004 -2804
rect 41404 -2806 42004 -2804
rect 77404 -2806 78004 -2804
rect 113404 -2806 114004 -2804
rect 149404 -2806 150004 -2804
rect 185404 -2806 186004 -2804
rect 221404 -2806 222004 -2804
rect 257404 -2806 258004 -2804
rect 293404 -2806 294004 -2804
rect 329404 -2806 330004 -2804
rect 365404 -2806 366004 -2804
rect 401404 -2806 402004 -2804
rect 437404 -2806 438004 -2804
rect 473404 -2806 474004 -2804
rect 509404 -2806 510004 -2804
rect 545404 -2806 546004 -2804
rect 581404 -2806 582004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 23404 -3144 24004 -3142
rect 59404 -3144 60004 -3142
rect 95404 -3144 96004 -3142
rect 131404 -3144 132004 -3142
rect 167404 -3144 168004 -3142
rect 203404 -3144 204004 -3142
rect 239404 -3144 240004 -3142
rect 275404 -3144 276004 -3142
rect 311404 -3144 312004 -3142
rect 347404 -3144 348004 -3142
rect 383404 -3144 384004 -3142
rect 419404 -3144 420004 -3142
rect 455404 -3144 456004 -3142
rect 491404 -3144 492004 -3142
rect 527404 -3144 528004 -3142
rect 563404 -3144 564004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3746 -4216 -3744
rect 23404 -3746 24004 -3744
rect 59404 -3746 60004 -3744
rect 95404 -3746 96004 -3744
rect 131404 -3746 132004 -3744
rect 167404 -3746 168004 -3744
rect 203404 -3746 204004 -3744
rect 239404 -3746 240004 -3744
rect 275404 -3746 276004 -3744
rect 311404 -3746 312004 -3744
rect 347404 -3746 348004 -3744
rect 383404 -3746 384004 -3744
rect 419404 -3746 420004 -3744
rect 455404 -3746 456004 -3744
rect 491404 -3746 492004 -3744
rect 527404 -3746 528004 -3744
rect 563404 -3746 564004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 9004 -4084 9604 -4082
rect 45004 -4084 45604 -4082
rect 81004 -4084 81604 -4082
rect 117004 -4084 117604 -4082
rect 153004 -4084 153604 -4082
rect 189004 -4084 189604 -4082
rect 225004 -4084 225604 -4082
rect 261004 -4084 261604 -4082
rect 297004 -4084 297604 -4082
rect 333004 -4084 333604 -4082
rect 369004 -4084 369604 -4082
rect 405004 -4084 405604 -4082
rect 441004 -4084 441604 -4082
rect 477004 -4084 477604 -4082
rect 513004 -4084 513604 -4082
rect 549004 -4084 549604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4686 -5156 -4684
rect 9004 -4686 9604 -4684
rect 45004 -4686 45604 -4684
rect 81004 -4686 81604 -4684
rect 117004 -4686 117604 -4684
rect 153004 -4686 153604 -4684
rect 189004 -4686 189604 -4684
rect 225004 -4686 225604 -4684
rect 261004 -4686 261604 -4684
rect 297004 -4686 297604 -4684
rect 333004 -4686 333604 -4684
rect 369004 -4686 369604 -4684
rect 405004 -4686 405604 -4684
rect 441004 -4686 441604 -4684
rect 477004 -4686 477604 -4684
rect 513004 -4686 513604 -4684
rect 549004 -4686 549604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 27004 -5024 27604 -5022
rect 63004 -5024 63604 -5022
rect 99004 -5024 99604 -5022
rect 135004 -5024 135604 -5022
rect 171004 -5024 171604 -5022
rect 207004 -5024 207604 -5022
rect 243004 -5024 243604 -5022
rect 279004 -5024 279604 -5022
rect 315004 -5024 315604 -5022
rect 351004 -5024 351604 -5022
rect 387004 -5024 387604 -5022
rect 423004 -5024 423604 -5022
rect 459004 -5024 459604 -5022
rect 495004 -5024 495604 -5022
rect 531004 -5024 531604 -5022
rect 567004 -5024 567604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5626 -6096 -5624
rect 27004 -5626 27604 -5624
rect 63004 -5626 63604 -5624
rect 99004 -5626 99604 -5624
rect 135004 -5626 135604 -5624
rect 171004 -5626 171604 -5624
rect 207004 -5626 207604 -5624
rect 243004 -5626 243604 -5624
rect 279004 -5626 279604 -5624
rect 315004 -5626 315604 -5624
rect 351004 -5626 351604 -5624
rect 387004 -5626 387604 -5624
rect 423004 -5626 423604 -5624
rect 459004 -5626 459604 -5624
rect 495004 -5626 495604 -5624
rect 531004 -5626 531604 -5624
rect 567004 -5626 567604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 12604 -5964 13204 -5962
rect 48604 -5964 49204 -5962
rect 84604 -5964 85204 -5962
rect 120604 -5964 121204 -5962
rect 156604 -5964 157204 -5962
rect 192604 -5964 193204 -5962
rect 228604 -5964 229204 -5962
rect 264604 -5964 265204 -5962
rect 300604 -5964 301204 -5962
rect 336604 -5964 337204 -5962
rect 372604 -5964 373204 -5962
rect 408604 -5964 409204 -5962
rect 444604 -5964 445204 -5962
rect 480604 -5964 481204 -5962
rect 516604 -5964 517204 -5962
rect 552604 -5964 553204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -6566 -7036 -6564
rect 12604 -6566 13204 -6564
rect 48604 -6566 49204 -6564
rect 84604 -6566 85204 -6564
rect 120604 -6566 121204 -6564
rect 156604 -6566 157204 -6564
rect 192604 -6566 193204 -6564
rect 228604 -6566 229204 -6564
rect 264604 -6566 265204 -6564
rect 300604 -6566 301204 -6564
rect 336604 -6566 337204 -6564
rect 372604 -6566 373204 -6564
rect 408604 -6566 409204 -6564
rect 444604 -6566 445204 -6564
rect 480604 -6566 481204 -6564
rect 516604 -6566 517204 -6564
rect 552604 -6566 553204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 30604 -6904 31204 -6902
rect 66604 -6904 67204 -6902
rect 102604 -6904 103204 -6902
rect 138604 -6904 139204 -6902
rect 174604 -6904 175204 -6902
rect 210604 -6904 211204 -6902
rect 246604 -6904 247204 -6902
rect 282604 -6904 283204 -6902
rect 318604 -6904 319204 -6902
rect 354604 -6904 355204 -6902
rect 390604 -6904 391204 -6902
rect 426604 -6904 427204 -6902
rect 462604 -6904 463204 -6902
rect 498604 -6904 499204 -6902
rect 534604 -6904 535204 -6902
rect 570604 -6904 571204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -7506 -7976 -7504
rect 30604 -7506 31204 -7504
rect 66604 -7506 67204 -7504
rect 102604 -7506 103204 -7504
rect 138604 -7506 139204 -7504
rect 174604 -7506 175204 -7504
rect 210604 -7506 211204 -7504
rect 246604 -7506 247204 -7504
rect 282604 -7506 283204 -7504
rect 318604 -7506 319204 -7504
rect 354604 -7506 355204 -7504
rect 390604 -7506 391204 -7504
rect 426604 -7506 427204 -7504
rect 462604 -7506 463204 -7504
rect 498604 -7506 499204 -7504
rect 534604 -7506 535204 -7504
rect 570604 -7506 571204 -7504
rect 591900 -7506 592500 -7504
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 696268 480 696508 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 636428 480 636668 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 576452 480 576692 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 516612 480 516852 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 456636 480 456876 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 681308 480 681548 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 621468 480 621708 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 561492 480 561732 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 501652 480 501892 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 441676 480 441916 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 396796 480 397036 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 351780 480 352020 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 306900 480 307140 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 262020 480 262260 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 217004 480 217244 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 172124 480 172364 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 127244 480 127484 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 82228 480 82468 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 37348 480 37588 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 651388 480 651628 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 591412 480 591652 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 531572 480 531812 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 471596 480 471836 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 411756 480 411996 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 366876 480 367116 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 321860 480 322100 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 276980 480 277220 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 231964 480 232204 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 187084 480 187324 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 142204 480 142444 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 97188 480 97428 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 52308 480 52548 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 7428 480 7668 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 666348 480 666588 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 606508 480 606748 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 546532 480 546772 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 486692 480 486932 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 426716 480 426956 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 381836 480 382076 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 336820 480 337060 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 291940 480 292180 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 247060 480 247300 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 202044 480 202284 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 157164 480 157404 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 112148 480 112388 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 67268 480 67508 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 22388 480 22628 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 400 nsew signal input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 401 nsew signal input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 402 nsew signal input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 403 nsew signal input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 404 nsew signal input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 405 nsew signal input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 406 nsew signal input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 407 nsew signal input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 408 nsew signal input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 409 nsew signal input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 410 nsew signal input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 411 nsew signal input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 412 nsew signal input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 413 nsew signal input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 414 nsew signal input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 415 nsew signal input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 416 nsew signal input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 417 nsew signal input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 418 nsew signal input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 419 nsew signal input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 420 nsew signal input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 421 nsew signal input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 422 nsew signal input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 423 nsew signal input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 424 nsew signal input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 425 nsew signal input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 426 nsew signal input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 427 nsew signal input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 429 nsew signal input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 430 nsew signal input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 431 nsew signal input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 432 nsew signal input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 433 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 434 nsew signal input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 435 nsew signal input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 436 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 437 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 438 nsew signal input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 439 nsew signal input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 440 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 441 nsew signal input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 442 nsew signal input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 443 nsew signal input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 444 nsew signal input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 445 nsew signal input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 446 nsew signal input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 447 nsew signal input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 448 nsew signal input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 449 nsew signal input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 450 nsew signal input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 451 nsew signal input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 452 nsew signal input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 453 nsew signal input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 454 nsew signal input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 455 nsew signal input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 456 nsew signal input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 457 nsew signal input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 458 nsew signal input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 459 nsew signal input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 460 nsew signal input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 461 nsew signal input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 462 nsew signal input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 463 nsew signal input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 464 nsew signal input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 465 nsew signal input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 466 nsew signal input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 467 nsew signal input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 468 nsew signal input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 469 nsew signal input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 470 nsew signal input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 471 nsew signal input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 472 nsew signal input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 473 nsew signal input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 474 nsew signal input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 475 nsew signal input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 476 nsew signal input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 477 nsew signal input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 478 nsew signal input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 479 nsew signal input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 480 nsew signal input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 481 nsew signal input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 482 nsew signal input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 483 nsew signal input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 484 nsew signal input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 485 nsew signal input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 486 nsew signal input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 487 nsew signal input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 488 nsew signal input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 489 nsew signal input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 490 nsew signal input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 491 nsew signal input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 492 nsew signal input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 493 nsew signal input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 494 nsew signal input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 495 nsew signal input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 496 nsew signal input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 497 nsew signal input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 498 nsew signal input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 499 nsew signal input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 500 nsew signal input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 501 nsew signal input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 502 nsew signal input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 503 nsew signal input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 504 nsew signal input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 505 nsew signal input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 506 nsew signal input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 507 nsew signal input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 508 nsew signal input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 509 nsew signal input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 510 nsew signal input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 511 nsew signal input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 512 nsew signal input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 513 nsew signal input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 514 nsew signal input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 515 nsew signal input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 516 nsew signal input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 517 nsew signal input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 518 nsew signal input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 519 nsew signal input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 520 nsew signal input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 521 nsew signal input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 522 nsew signal input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 523 nsew signal input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 524 nsew signal input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 525 nsew signal input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 526 nsew signal input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 527 nsew signal input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 529 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 530 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 531 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 532 nsew signal input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 533 nsew signal input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 534 nsew signal input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 535 nsew signal input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 536 nsew signal input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 537 nsew signal input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 538 nsew signal input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 539 nsew signal input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 540 nsew signal input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 541 nsew signal input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 542 nsew signal input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 543 nsew signal input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 544 nsew signal input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 545 nsew signal input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 546 nsew signal input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 547 nsew signal input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 548 nsew signal input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 549 nsew signal input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 550 nsew signal input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 551 nsew signal input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 552 nsew signal input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 553 nsew signal input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 554 nsew signal input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 555 nsew signal input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 556 nsew signal input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 557 nsew signal input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 558 nsew signal input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 559 nsew signal input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 560 nsew signal input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 561 nsew signal input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 562 nsew signal input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 563 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 564 nsew signal input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 565 nsew signal input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 566 nsew signal input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 567 nsew signal input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 568 nsew signal input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 569 nsew signal input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 570 nsew signal input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 571 nsew signal input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 572 nsew signal input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 573 nsew signal input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 574 nsew signal input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 575 nsew signal input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 576 nsew signal input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 577 nsew signal input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 578 nsew signal input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 579 nsew signal input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 580 nsew signal input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 581 nsew signal input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 582 nsew signal input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 583 nsew signal input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 584 nsew signal input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 585 nsew signal input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 586 nsew signal input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 587 nsew signal input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 588 nsew signal input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 589 nsew signal input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 590 nsew signal input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 591 nsew signal input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 592 nsew signal input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 593 nsew signal input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 594 nsew signal input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 595 nsew signal input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 596 nsew signal input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 597 nsew signal output
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 598 nsew signal output
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 599 nsew signal output
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 600 nsew signal output
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 601 nsew signal output
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 602 nsew signal output
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 603 nsew signal output
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 604 nsew signal output
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 605 nsew signal output
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 606 nsew signal output
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 607 nsew signal output
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 608 nsew signal output
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 609 nsew signal output
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 610 nsew signal output
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 611 nsew signal output
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 612 nsew signal output
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 613 nsew signal output
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 614 nsew signal output
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 615 nsew signal output
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 616 nsew signal output
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 617 nsew signal output
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 618 nsew signal output
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 619 nsew signal output
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 620 nsew signal output
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 621 nsew signal output
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 622 nsew signal output
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 623 nsew signal output
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 624 nsew signal output
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 625 nsew signal output
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 626 nsew signal output
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 627 nsew signal output
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 628 nsew signal output
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 629 nsew signal input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 630 nsew signal input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 631 nsew signal input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 632 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 633 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 634 nsew signal input
rlabel metal4 s 577804 -1864 578404 705800 6 vccd1
port 635 nsew power bidirectional
rlabel metal4 s 541804 -1864 542404 705800 6 vccd1
port 636 nsew power bidirectional
rlabel metal4 s 505804 613152 506404 705800 6 vccd1
port 637 nsew power bidirectional
rlabel metal4 s 469804 613152 470404 705800 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 433804 -1864 434404 705800 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 397804 -1864 398404 705800 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 361804 613152 362404 705800 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 325804 613152 326404 705800 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s 289804 -1864 290404 705800 6 vccd1
port 643 nsew power bidirectional
rlabel metal4 s 253804 613152 254404 705800 6 vccd1
port 644 nsew power bidirectional
rlabel metal4 s 217804 613152 218404 705800 6 vccd1
port 645 nsew power bidirectional
rlabel metal4 s 181804 -1864 182404 705800 6 vccd1
port 646 nsew power bidirectional
rlabel metal4 s 145804 -1864 146404 705800 6 vccd1
port 647 nsew power bidirectional
rlabel metal4 s 109804 613152 110404 705800 6 vccd1
port 648 nsew power bidirectional
rlabel metal4 s 73804 613152 74404 705800 6 vccd1
port 649 nsew power bidirectional
rlabel metal4 s 37804 -1864 38404 705800 6 vccd1
port 650 nsew power bidirectional
rlabel metal4 s 1804 -1864 2404 705800 6 vccd1
port 651 nsew power bidirectional
rlabel metal4 s 585320 -924 585920 704860 6 vccd1
port 652 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1
port 653 nsew power bidirectional
rlabel metal4 s 505804 460352 506404 549248 6 vccd1
port 654 nsew power bidirectional
rlabel metal4 s 469804 460352 470404 549248 6 vccd1
port 655 nsew power bidirectional
rlabel metal4 s 361804 460352 362404 549248 6 vccd1
port 656 nsew power bidirectional
rlabel metal4 s 325804 460352 326404 549248 6 vccd1
port 657 nsew power bidirectional
rlabel metal4 s 253804 460352 254404 549248 6 vccd1
port 658 nsew power bidirectional
rlabel metal4 s 217804 460352 218404 549248 6 vccd1
port 659 nsew power bidirectional
rlabel metal4 s 109804 460352 110404 549248 6 vccd1
port 660 nsew power bidirectional
rlabel metal4 s 73804 460352 74404 549248 6 vccd1
port 661 nsew power bidirectional
rlabel metal4 s 505804 307552 506404 396448 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 469804 307552 470404 396448 6 vccd1
port 663 nsew power bidirectional
rlabel metal4 s 361804 307552 362404 396448 6 vccd1
port 664 nsew power bidirectional
rlabel metal4 s 325804 307552 326404 396448 6 vccd1
port 665 nsew power bidirectional
rlabel metal4 s 253804 307552 254404 396448 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 217804 307552 218404 396448 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 109804 307552 110404 396448 6 vccd1
port 668 nsew power bidirectional
rlabel metal4 s 73804 307552 74404 396448 6 vccd1
port 669 nsew power bidirectional
rlabel metal4 s 505804 154752 506404 243648 6 vccd1
port 670 nsew power bidirectional
rlabel metal4 s 469804 154752 470404 243648 6 vccd1
port 671 nsew power bidirectional
rlabel metal4 s 361804 154752 362404 243648 6 vccd1
port 672 nsew power bidirectional
rlabel metal4 s 325804 154752 326404 243648 6 vccd1
port 673 nsew power bidirectional
rlabel metal4 s 253804 154752 254404 243648 6 vccd1
port 674 nsew power bidirectional
rlabel metal4 s 217804 154752 218404 243648 6 vccd1
port 675 nsew power bidirectional
rlabel metal4 s 109804 154752 110404 243648 6 vccd1
port 676 nsew power bidirectional
rlabel metal4 s 73804 154752 74404 243648 6 vccd1
port 677 nsew power bidirectional
rlabel metal4 s 505804 -1864 506404 90848 6 vccd1
port 678 nsew power bidirectional
rlabel metal4 s 469804 -1864 470404 90848 6 vccd1
port 679 nsew power bidirectional
rlabel metal4 s 361804 -1864 362404 90848 6 vccd1
port 680 nsew power bidirectional
rlabel metal4 s 325804 -1864 326404 90848 6 vccd1
port 681 nsew power bidirectional
rlabel metal4 s 253804 -1864 254404 90848 6 vccd1
port 682 nsew power bidirectional
rlabel metal4 s 217804 -1864 218404 90848 6 vccd1
port 683 nsew power bidirectional
rlabel metal4 s 109804 -1864 110404 90848 6 vccd1
port 684 nsew power bidirectional
rlabel metal4 s 73804 -1864 74404 90848 6 vccd1
port 685 nsew power bidirectional
rlabel metal5 s -1996 704260 585920 704860 6 vccd1
port 686 nsew power bidirectional
rlabel metal5 s -2936 686828 586860 687428 6 vccd1
port 687 nsew power bidirectional
rlabel metal5 s -2936 650828 586860 651428 6 vccd1
port 688 nsew power bidirectional
rlabel metal5 s -2936 614828 586860 615428 6 vccd1
port 689 nsew power bidirectional
rlabel metal5 s -2936 578828 586860 579428 6 vccd1
port 690 nsew power bidirectional
rlabel metal5 s -2936 542828 586860 543428 6 vccd1
port 691 nsew power bidirectional
rlabel metal5 s -2936 506828 586860 507428 6 vccd1
port 692 nsew power bidirectional
rlabel metal5 s -2936 470828 586860 471428 6 vccd1
port 693 nsew power bidirectional
rlabel metal5 s -2936 434828 586860 435428 6 vccd1
port 694 nsew power bidirectional
rlabel metal5 s -2936 398828 586860 399428 6 vccd1
port 695 nsew power bidirectional
rlabel metal5 s -2936 362828 586860 363428 6 vccd1
port 696 nsew power bidirectional
rlabel metal5 s -2936 326828 586860 327428 6 vccd1
port 697 nsew power bidirectional
rlabel metal5 s -2936 290828 586860 291428 6 vccd1
port 698 nsew power bidirectional
rlabel metal5 s -2936 254828 586860 255428 6 vccd1
port 699 nsew power bidirectional
rlabel metal5 s -2936 218828 586860 219428 6 vccd1
port 700 nsew power bidirectional
rlabel metal5 s -2936 182828 586860 183428 6 vccd1
port 701 nsew power bidirectional
rlabel metal5 s -2936 146828 586860 147428 6 vccd1
port 702 nsew power bidirectional
rlabel metal5 s -2936 110828 586860 111428 6 vccd1
port 703 nsew power bidirectional
rlabel metal5 s -2936 74828 586860 75428 6 vccd1
port 704 nsew power bidirectional
rlabel metal5 s -2936 38828 586860 39428 6 vccd1
port 705 nsew power bidirectional
rlabel metal5 s -2936 2828 586860 3428 6 vccd1
port 706 nsew power bidirectional
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 707 nsew power bidirectional
rlabel metal4 s 586260 -1864 586860 705800 6 vssd1
port 708 nsew ground bidirectional
rlabel metal4 s 559804 -1864 560404 705800 6 vssd1
port 709 nsew ground bidirectional
rlabel metal4 s 523804 -1864 524404 705800 6 vssd1
port 710 nsew ground bidirectional
rlabel metal4 s 487804 613152 488404 705800 6 vssd1
port 711 nsew ground bidirectional
rlabel metal4 s 451804 -1864 452404 705800 6 vssd1
port 712 nsew ground bidirectional
rlabel metal4 s 415804 -1864 416404 705800 6 vssd1
port 713 nsew ground bidirectional
rlabel metal4 s 379804 613152 380404 705800 6 vssd1
port 714 nsew ground bidirectional
rlabel metal4 s 343804 613152 344404 705800 6 vssd1
port 715 nsew ground bidirectional
rlabel metal4 s 307804 -1864 308404 705800 6 vssd1
port 716 nsew ground bidirectional
rlabel metal4 s 271804 -1864 272404 705800 6 vssd1
port 717 nsew ground bidirectional
rlabel metal4 s 235804 613152 236404 705800 6 vssd1
port 718 nsew ground bidirectional
rlabel metal4 s 199804 613152 200404 705800 6 vssd1
port 719 nsew ground bidirectional
rlabel metal4 s 163804 -1864 164404 705800 6 vssd1
port 720 nsew ground bidirectional
rlabel metal4 s 127804 613152 128404 705800 6 vssd1
port 721 nsew ground bidirectional
rlabel metal4 s 91804 613152 92404 705800 6 vssd1
port 722 nsew ground bidirectional
rlabel metal4 s 55804 -1864 56404 705800 6 vssd1
port 723 nsew ground bidirectional
rlabel metal4 s 19804 -1864 20404 705800 6 vssd1
port 724 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1
port 725 nsew ground bidirectional
rlabel metal4 s 487804 460352 488404 549248 6 vssd1
port 726 nsew ground bidirectional
rlabel metal4 s 379804 460352 380404 549248 6 vssd1
port 727 nsew ground bidirectional
rlabel metal4 s 343804 460352 344404 549248 6 vssd1
port 728 nsew ground bidirectional
rlabel metal4 s 235804 460352 236404 549248 6 vssd1
port 729 nsew ground bidirectional
rlabel metal4 s 199804 460352 200404 549248 6 vssd1
port 730 nsew ground bidirectional
rlabel metal4 s 127804 460352 128404 549248 6 vssd1
port 731 nsew ground bidirectional
rlabel metal4 s 91804 460352 92404 549248 6 vssd1
port 732 nsew ground bidirectional
rlabel metal4 s 487804 307552 488404 396448 6 vssd1
port 733 nsew ground bidirectional
rlabel metal4 s 379804 307552 380404 396448 6 vssd1
port 734 nsew ground bidirectional
rlabel metal4 s 343804 307552 344404 396448 6 vssd1
port 735 nsew ground bidirectional
rlabel metal4 s 235804 307552 236404 396448 6 vssd1
port 736 nsew ground bidirectional
rlabel metal4 s 199804 307552 200404 396448 6 vssd1
port 737 nsew ground bidirectional
rlabel metal4 s 127804 307552 128404 396448 6 vssd1
port 738 nsew ground bidirectional
rlabel metal4 s 91804 307552 92404 396448 6 vssd1
port 739 nsew ground bidirectional
rlabel metal4 s 487804 154752 488404 243648 6 vssd1
port 740 nsew ground bidirectional
rlabel metal4 s 379804 154752 380404 243648 6 vssd1
port 741 nsew ground bidirectional
rlabel metal4 s 343804 154752 344404 243648 6 vssd1
port 742 nsew ground bidirectional
rlabel metal4 s 235804 154752 236404 243648 6 vssd1
port 743 nsew ground bidirectional
rlabel metal4 s 199804 154752 200404 243648 6 vssd1
port 744 nsew ground bidirectional
rlabel metal4 s 127804 154752 128404 243648 6 vssd1
port 745 nsew ground bidirectional
rlabel metal4 s 91804 154752 92404 243648 6 vssd1
port 746 nsew ground bidirectional
rlabel metal4 s 487804 -1864 488404 90848 6 vssd1
port 747 nsew ground bidirectional
rlabel metal4 s 379804 -1864 380404 90848 6 vssd1
port 748 nsew ground bidirectional
rlabel metal4 s 343804 -1864 344404 90848 6 vssd1
port 749 nsew ground bidirectional
rlabel metal4 s 235804 -1864 236404 90848 6 vssd1
port 750 nsew ground bidirectional
rlabel metal4 s 199804 -1864 200404 90848 6 vssd1
port 751 nsew ground bidirectional
rlabel metal4 s 127804 -1864 128404 90848 6 vssd1
port 752 nsew ground bidirectional
rlabel metal4 s 91804 -1864 92404 90848 6 vssd1
port 753 nsew ground bidirectional
rlabel metal5 s -2936 705200 586860 705800 6 vssd1
port 754 nsew ground bidirectional
rlabel metal5 s -2936 668828 586860 669428 6 vssd1
port 755 nsew ground bidirectional
rlabel metal5 s -2936 632828 586860 633428 6 vssd1
port 756 nsew ground bidirectional
rlabel metal5 s -2936 596828 586860 597428 6 vssd1
port 757 nsew ground bidirectional
rlabel metal5 s -2936 560828 586860 561428 6 vssd1
port 758 nsew ground bidirectional
rlabel metal5 s -2936 524828 586860 525428 6 vssd1
port 759 nsew ground bidirectional
rlabel metal5 s -2936 488828 586860 489428 6 vssd1
port 760 nsew ground bidirectional
rlabel metal5 s -2936 452828 586860 453428 6 vssd1
port 761 nsew ground bidirectional
rlabel metal5 s -2936 416828 586860 417428 6 vssd1
port 762 nsew ground bidirectional
rlabel metal5 s -2936 380828 586860 381428 6 vssd1
port 763 nsew ground bidirectional
rlabel metal5 s -2936 344828 586860 345428 6 vssd1
port 764 nsew ground bidirectional
rlabel metal5 s -2936 308828 586860 309428 6 vssd1
port 765 nsew ground bidirectional
rlabel metal5 s -2936 272828 586860 273428 6 vssd1
port 766 nsew ground bidirectional
rlabel metal5 s -2936 236828 586860 237428 6 vssd1
port 767 nsew ground bidirectional
rlabel metal5 s -2936 200828 586860 201428 6 vssd1
port 768 nsew ground bidirectional
rlabel metal5 s -2936 164828 586860 165428 6 vssd1
port 769 nsew ground bidirectional
rlabel metal5 s -2936 128828 586860 129428 6 vssd1
port 770 nsew ground bidirectional
rlabel metal5 s -2936 92828 586860 93428 6 vssd1
port 771 nsew ground bidirectional
rlabel metal5 s -2936 56828 586860 57428 6 vssd1
port 772 nsew ground bidirectional
rlabel metal5 s -2936 20828 586860 21428 6 vssd1
port 773 nsew ground bidirectional
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 774 nsew ground bidirectional
rlabel metal4 s 581404 -3744 582004 707680 6 vccd2
port 775 nsew power bidirectional
rlabel metal4 s 545404 -3744 546004 707680 6 vccd2
port 776 nsew power bidirectional
rlabel metal4 s 509404 613200 510004 707680 6 vccd2
port 777 nsew power bidirectional
rlabel metal4 s 473404 613200 474004 707680 6 vccd2
port 778 nsew power bidirectional
rlabel metal4 s 437404 -3744 438004 707680 6 vccd2
port 779 nsew power bidirectional
rlabel metal4 s 401404 -3744 402004 707680 6 vccd2
port 780 nsew power bidirectional
rlabel metal4 s 365404 613200 366004 707680 6 vccd2
port 781 nsew power bidirectional
rlabel metal4 s 329404 613200 330004 707680 6 vccd2
port 782 nsew power bidirectional
rlabel metal4 s 293404 -3744 294004 707680 6 vccd2
port 783 nsew power bidirectional
rlabel metal4 s 257404 613200 258004 707680 6 vccd2
port 784 nsew power bidirectional
rlabel metal4 s 221404 613200 222004 707680 6 vccd2
port 785 nsew power bidirectional
rlabel metal4 s 185404 -3744 186004 707680 6 vccd2
port 786 nsew power bidirectional
rlabel metal4 s 149404 -3744 150004 707680 6 vccd2
port 787 nsew power bidirectional
rlabel metal4 s 113404 613200 114004 707680 6 vccd2
port 788 nsew power bidirectional
rlabel metal4 s 77404 613200 78004 707680 6 vccd2
port 789 nsew power bidirectional
rlabel metal4 s 41404 -3744 42004 707680 6 vccd2
port 790 nsew power bidirectional
rlabel metal4 s 5404 -3744 6004 707680 6 vccd2
port 791 nsew power bidirectional
rlabel metal4 s 587200 -2804 587800 706740 6 vccd2
port 792 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2
port 793 nsew power bidirectional
rlabel metal4 s 509404 460400 510004 549200 6 vccd2
port 794 nsew power bidirectional
rlabel metal4 s 473404 460400 474004 549200 6 vccd2
port 795 nsew power bidirectional
rlabel metal4 s 365404 460400 366004 549200 6 vccd2
port 796 nsew power bidirectional
rlabel metal4 s 329404 460400 330004 549200 6 vccd2
port 797 nsew power bidirectional
rlabel metal4 s 257404 460400 258004 549200 6 vccd2
port 798 nsew power bidirectional
rlabel metal4 s 221404 460400 222004 549200 6 vccd2
port 799 nsew power bidirectional
rlabel metal4 s 113404 460400 114004 549200 6 vccd2
port 800 nsew power bidirectional
rlabel metal4 s 77404 460400 78004 549200 6 vccd2
port 801 nsew power bidirectional
rlabel metal4 s 509404 307600 510004 396400 6 vccd2
port 802 nsew power bidirectional
rlabel metal4 s 473404 307600 474004 396400 6 vccd2
port 803 nsew power bidirectional
rlabel metal4 s 365404 307600 366004 396400 6 vccd2
port 804 nsew power bidirectional
rlabel metal4 s 329404 307600 330004 396400 6 vccd2
port 805 nsew power bidirectional
rlabel metal4 s 257404 307600 258004 396400 6 vccd2
port 806 nsew power bidirectional
rlabel metal4 s 221404 307600 222004 396400 6 vccd2
port 807 nsew power bidirectional
rlabel metal4 s 113404 307600 114004 396400 6 vccd2
port 808 nsew power bidirectional
rlabel metal4 s 77404 307600 78004 396400 6 vccd2
port 809 nsew power bidirectional
rlabel metal4 s 509404 154800 510004 243600 6 vccd2
port 810 nsew power bidirectional
rlabel metal4 s 473404 154800 474004 243600 6 vccd2
port 811 nsew power bidirectional
rlabel metal4 s 365404 154800 366004 243600 6 vccd2
port 812 nsew power bidirectional
rlabel metal4 s 329404 154800 330004 243600 6 vccd2
port 813 nsew power bidirectional
rlabel metal4 s 257404 154800 258004 243600 6 vccd2
port 814 nsew power bidirectional
rlabel metal4 s 221404 154800 222004 243600 6 vccd2
port 815 nsew power bidirectional
rlabel metal4 s 113404 154800 114004 243600 6 vccd2
port 816 nsew power bidirectional
rlabel metal4 s 77404 154800 78004 243600 6 vccd2
port 817 nsew power bidirectional
rlabel metal4 s 509404 -3744 510004 90800 6 vccd2
port 818 nsew power bidirectional
rlabel metal4 s 473404 -3744 474004 90800 6 vccd2
port 819 nsew power bidirectional
rlabel metal4 s 365404 -3744 366004 90800 6 vccd2
port 820 nsew power bidirectional
rlabel metal4 s 329404 -3744 330004 90800 6 vccd2
port 821 nsew power bidirectional
rlabel metal4 s 257404 -3744 258004 90800 6 vccd2
port 822 nsew power bidirectional
rlabel metal4 s 221404 -3744 222004 90800 6 vccd2
port 823 nsew power bidirectional
rlabel metal4 s 113404 -3744 114004 90800 6 vccd2
port 824 nsew power bidirectional
rlabel metal4 s 77404 -3744 78004 90800 6 vccd2
port 825 nsew power bidirectional
rlabel metal5 s -3876 706140 587800 706740 6 vccd2
port 826 nsew power bidirectional
rlabel metal5 s -4816 690476 588740 691076 6 vccd2
port 827 nsew power bidirectional
rlabel metal5 s -4816 654476 588740 655076 6 vccd2
port 828 nsew power bidirectional
rlabel metal5 s -4816 618476 588740 619076 6 vccd2
port 829 nsew power bidirectional
rlabel metal5 s -4816 582476 588740 583076 6 vccd2
port 830 nsew power bidirectional
rlabel metal5 s -4816 546476 588740 547076 6 vccd2
port 831 nsew power bidirectional
rlabel metal5 s -4816 510476 588740 511076 6 vccd2
port 832 nsew power bidirectional
rlabel metal5 s -4816 474476 588740 475076 6 vccd2
port 833 nsew power bidirectional
rlabel metal5 s -4816 438476 588740 439076 6 vccd2
port 834 nsew power bidirectional
rlabel metal5 s -4816 402476 588740 403076 6 vccd2
port 835 nsew power bidirectional
rlabel metal5 s -4816 366476 588740 367076 6 vccd2
port 836 nsew power bidirectional
rlabel metal5 s -4816 330476 588740 331076 6 vccd2
port 837 nsew power bidirectional
rlabel metal5 s -4816 294476 588740 295076 6 vccd2
port 838 nsew power bidirectional
rlabel metal5 s -4816 258476 588740 259076 6 vccd2
port 839 nsew power bidirectional
rlabel metal5 s -4816 222476 588740 223076 6 vccd2
port 840 nsew power bidirectional
rlabel metal5 s -4816 186476 588740 187076 6 vccd2
port 841 nsew power bidirectional
rlabel metal5 s -4816 150476 588740 151076 6 vccd2
port 842 nsew power bidirectional
rlabel metal5 s -4816 114476 588740 115076 6 vccd2
port 843 nsew power bidirectional
rlabel metal5 s -4816 78476 588740 79076 6 vccd2
port 844 nsew power bidirectional
rlabel metal5 s -4816 42476 588740 43076 6 vccd2
port 845 nsew power bidirectional
rlabel metal5 s -4816 6476 588740 7076 6 vccd2
port 846 nsew power bidirectional
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 847 nsew power bidirectional
rlabel metal4 s 588140 -3744 588740 707680 6 vssd2
port 848 nsew ground bidirectional
rlabel metal4 s 563404 -3744 564004 707680 6 vssd2
port 849 nsew ground bidirectional
rlabel metal4 s 527404 -3744 528004 707680 6 vssd2
port 850 nsew ground bidirectional
rlabel metal4 s 491404 613200 492004 707680 6 vssd2
port 851 nsew ground bidirectional
rlabel metal4 s 455404 613200 456004 707680 6 vssd2
port 852 nsew ground bidirectional
rlabel metal4 s 419404 -3744 420004 707680 6 vssd2
port 853 nsew ground bidirectional
rlabel metal4 s 383404 613200 384004 707680 6 vssd2
port 854 nsew ground bidirectional
rlabel metal4 s 347404 613200 348004 707680 6 vssd2
port 855 nsew ground bidirectional
rlabel metal4 s 311404 -3744 312004 707680 6 vssd2
port 856 nsew ground bidirectional
rlabel metal4 s 275404 -3744 276004 707680 6 vssd2
port 857 nsew ground bidirectional
rlabel metal4 s 239404 613200 240004 707680 6 vssd2
port 858 nsew ground bidirectional
rlabel metal4 s 203404 613200 204004 707680 6 vssd2
port 859 nsew ground bidirectional
rlabel metal4 s 167404 -3744 168004 707680 6 vssd2
port 860 nsew ground bidirectional
rlabel metal4 s 131404 -3744 132004 707680 6 vssd2
port 861 nsew ground bidirectional
rlabel metal4 s 95404 613200 96004 707680 6 vssd2
port 862 nsew ground bidirectional
rlabel metal4 s 59404 -3744 60004 707680 6 vssd2
port 863 nsew ground bidirectional
rlabel metal4 s 23404 -3744 24004 707680 6 vssd2
port 864 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2
port 865 nsew ground bidirectional
rlabel metal4 s 491404 460400 492004 549200 6 vssd2
port 866 nsew ground bidirectional
rlabel metal4 s 455404 460400 456004 549200 6 vssd2
port 867 nsew ground bidirectional
rlabel metal4 s 383404 460400 384004 549200 6 vssd2
port 868 nsew ground bidirectional
rlabel metal4 s 347404 460400 348004 549200 6 vssd2
port 869 nsew ground bidirectional
rlabel metal4 s 239404 460400 240004 549200 6 vssd2
port 870 nsew ground bidirectional
rlabel metal4 s 203404 460400 204004 549200 6 vssd2
port 871 nsew ground bidirectional
rlabel metal4 s 95404 460400 96004 549200 6 vssd2
port 872 nsew ground bidirectional
rlabel metal4 s 491404 307600 492004 396400 6 vssd2
port 873 nsew ground bidirectional
rlabel metal4 s 455404 307600 456004 396400 6 vssd2
port 874 nsew ground bidirectional
rlabel metal4 s 383404 307600 384004 396400 6 vssd2
port 875 nsew ground bidirectional
rlabel metal4 s 347404 307600 348004 396400 6 vssd2
port 876 nsew ground bidirectional
rlabel metal4 s 239404 307600 240004 396400 6 vssd2
port 877 nsew ground bidirectional
rlabel metal4 s 203404 307600 204004 396400 6 vssd2
port 878 nsew ground bidirectional
rlabel metal4 s 95404 307600 96004 396400 6 vssd2
port 879 nsew ground bidirectional
rlabel metal4 s 491404 154800 492004 243600 6 vssd2
port 880 nsew ground bidirectional
rlabel metal4 s 455404 154800 456004 243600 6 vssd2
port 881 nsew ground bidirectional
rlabel metal4 s 383404 154800 384004 243600 6 vssd2
port 882 nsew ground bidirectional
rlabel metal4 s 347404 154800 348004 243600 6 vssd2
port 883 nsew ground bidirectional
rlabel metal4 s 239404 154800 240004 243600 6 vssd2
port 884 nsew ground bidirectional
rlabel metal4 s 203404 154800 204004 243600 6 vssd2
port 885 nsew ground bidirectional
rlabel metal4 s 95404 154800 96004 243600 6 vssd2
port 886 nsew ground bidirectional
rlabel metal4 s 491404 -3744 492004 90800 6 vssd2
port 887 nsew ground bidirectional
rlabel metal4 s 455404 -3744 456004 90800 6 vssd2
port 888 nsew ground bidirectional
rlabel metal4 s 383404 -3744 384004 90800 6 vssd2
port 889 nsew ground bidirectional
rlabel metal4 s 347404 -3744 348004 90800 6 vssd2
port 890 nsew ground bidirectional
rlabel metal4 s 239404 -3744 240004 90800 6 vssd2
port 891 nsew ground bidirectional
rlabel metal4 s 203404 -3744 204004 90800 6 vssd2
port 892 nsew ground bidirectional
rlabel metal4 s 95404 -3744 96004 90800 6 vssd2
port 893 nsew ground bidirectional
rlabel metal5 s -4816 707080 588740 707680 6 vssd2
port 894 nsew ground bidirectional
rlabel metal5 s -4816 672476 588740 673076 6 vssd2
port 895 nsew ground bidirectional
rlabel metal5 s -4816 636476 588740 637076 6 vssd2
port 896 nsew ground bidirectional
rlabel metal5 s -4816 600476 588740 601076 6 vssd2
port 897 nsew ground bidirectional
rlabel metal5 s -4816 564476 588740 565076 6 vssd2
port 898 nsew ground bidirectional
rlabel metal5 s -4816 528476 588740 529076 6 vssd2
port 899 nsew ground bidirectional
rlabel metal5 s -4816 492476 588740 493076 6 vssd2
port 900 nsew ground bidirectional
rlabel metal5 s -4816 456476 588740 457076 6 vssd2
port 901 nsew ground bidirectional
rlabel metal5 s -4816 420476 588740 421076 6 vssd2
port 902 nsew ground bidirectional
rlabel metal5 s -4816 384476 588740 385076 6 vssd2
port 903 nsew ground bidirectional
rlabel metal5 s -4816 348476 588740 349076 6 vssd2
port 904 nsew ground bidirectional
rlabel metal5 s -4816 312476 588740 313076 6 vssd2
port 905 nsew ground bidirectional
rlabel metal5 s -4816 276476 588740 277076 6 vssd2
port 906 nsew ground bidirectional
rlabel metal5 s -4816 240476 588740 241076 6 vssd2
port 907 nsew ground bidirectional
rlabel metal5 s -4816 204476 588740 205076 6 vssd2
port 908 nsew ground bidirectional
rlabel metal5 s -4816 168476 588740 169076 6 vssd2
port 909 nsew ground bidirectional
rlabel metal5 s -4816 132476 588740 133076 6 vssd2
port 910 nsew ground bidirectional
rlabel metal5 s -4816 96476 588740 97076 6 vssd2
port 911 nsew ground bidirectional
rlabel metal5 s -4816 60476 588740 61076 6 vssd2
port 912 nsew ground bidirectional
rlabel metal5 s -4816 24476 588740 25076 6 vssd2
port 913 nsew ground bidirectional
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 914 nsew ground bidirectional
rlabel metal4 s 549004 -5624 549604 709560 6 vdda1
port 915 nsew power bidirectional
rlabel metal4 s 513004 613200 513604 709560 6 vdda1
port 916 nsew power bidirectional
rlabel metal4 s 477004 613200 477604 709560 6 vdda1
port 917 nsew power bidirectional
rlabel metal4 s 441004 -5624 441604 709560 6 vdda1
port 918 nsew power bidirectional
rlabel metal4 s 405004 -5624 405604 709560 6 vdda1
port 919 nsew power bidirectional
rlabel metal4 s 369004 613200 369604 709560 6 vdda1
port 920 nsew power bidirectional
rlabel metal4 s 333004 613200 333604 709560 6 vdda1
port 921 nsew power bidirectional
rlabel metal4 s 297004 -5624 297604 709560 6 vdda1
port 922 nsew power bidirectional
rlabel metal4 s 261004 -5624 261604 709560 6 vdda1
port 923 nsew power bidirectional
rlabel metal4 s 225004 613200 225604 709560 6 vdda1
port 924 nsew power bidirectional
rlabel metal4 s 189004 -5624 189604 709560 6 vdda1
port 925 nsew power bidirectional
rlabel metal4 s 153004 -5624 153604 709560 6 vdda1
port 926 nsew power bidirectional
rlabel metal4 s 117004 613200 117604 709560 6 vdda1
port 927 nsew power bidirectional
rlabel metal4 s 81004 613200 81604 709560 6 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 45004 -5624 45604 709560 6 vdda1
port 929 nsew power bidirectional
rlabel metal4 s 9004 -5624 9604 709560 6 vdda1
port 930 nsew power bidirectional
rlabel metal4 s 589080 -4684 589680 708620 6 vdda1
port 931 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1
port 932 nsew power bidirectional
rlabel metal4 s 513004 460400 513604 549200 6 vdda1
port 933 nsew power bidirectional
rlabel metal4 s 477004 460400 477604 549200 6 vdda1
port 934 nsew power bidirectional
rlabel metal4 s 369004 460400 369604 549200 6 vdda1
port 935 nsew power bidirectional
rlabel metal4 s 333004 460400 333604 549200 6 vdda1
port 936 nsew power bidirectional
rlabel metal4 s 225004 460400 225604 549200 6 vdda1
port 937 nsew power bidirectional
rlabel metal4 s 117004 460400 117604 549200 6 vdda1
port 938 nsew power bidirectional
rlabel metal4 s 81004 460400 81604 549200 6 vdda1
port 939 nsew power bidirectional
rlabel metal4 s 513004 307600 513604 396400 6 vdda1
port 940 nsew power bidirectional
rlabel metal4 s 477004 307600 477604 396400 6 vdda1
port 941 nsew power bidirectional
rlabel metal4 s 369004 307600 369604 396400 6 vdda1
port 942 nsew power bidirectional
rlabel metal4 s 333004 307600 333604 396400 6 vdda1
port 943 nsew power bidirectional
rlabel metal4 s 225004 307600 225604 396400 6 vdda1
port 944 nsew power bidirectional
rlabel metal4 s 117004 307600 117604 396400 6 vdda1
port 945 nsew power bidirectional
rlabel metal4 s 81004 307600 81604 396400 6 vdda1
port 946 nsew power bidirectional
rlabel metal4 s 513004 154800 513604 243600 6 vdda1
port 947 nsew power bidirectional
rlabel metal4 s 477004 154800 477604 243600 6 vdda1
port 948 nsew power bidirectional
rlabel metal4 s 369004 154800 369604 243600 6 vdda1
port 949 nsew power bidirectional
rlabel metal4 s 333004 154800 333604 243600 6 vdda1
port 950 nsew power bidirectional
rlabel metal4 s 225004 154800 225604 243600 6 vdda1
port 951 nsew power bidirectional
rlabel metal4 s 117004 154800 117604 243600 6 vdda1
port 952 nsew power bidirectional
rlabel metal4 s 81004 154800 81604 243600 6 vdda1
port 953 nsew power bidirectional
rlabel metal4 s 513004 -5624 513604 90800 6 vdda1
port 954 nsew power bidirectional
rlabel metal4 s 477004 -5624 477604 90800 6 vdda1
port 955 nsew power bidirectional
rlabel metal4 s 369004 -5624 369604 90800 6 vdda1
port 956 nsew power bidirectional
rlabel metal4 s 333004 -5624 333604 90800 6 vdda1
port 957 nsew power bidirectional
rlabel metal4 s 225004 -5624 225604 90800 6 vdda1
port 958 nsew power bidirectional
rlabel metal4 s 117004 -5624 117604 90800 6 vdda1
port 959 nsew power bidirectional
rlabel metal4 s 81004 -5624 81604 90800 6 vdda1
port 960 nsew power bidirectional
rlabel metal5 s -5756 708020 589680 708620 6 vdda1
port 961 nsew power bidirectional
rlabel metal5 s -6696 694076 590620 694676 6 vdda1
port 962 nsew power bidirectional
rlabel metal5 s -6696 658076 590620 658676 6 vdda1
port 963 nsew power bidirectional
rlabel metal5 s -6696 622076 590620 622676 6 vdda1
port 964 nsew power bidirectional
rlabel metal5 s -6696 586076 590620 586676 6 vdda1
port 965 nsew power bidirectional
rlabel metal5 s -6696 550076 590620 550676 6 vdda1
port 966 nsew power bidirectional
rlabel metal5 s -6696 514076 590620 514676 6 vdda1
port 967 nsew power bidirectional
rlabel metal5 s -6696 478076 590620 478676 6 vdda1
port 968 nsew power bidirectional
rlabel metal5 s -6696 442076 590620 442676 6 vdda1
port 969 nsew power bidirectional
rlabel metal5 s -6696 406076 590620 406676 6 vdda1
port 970 nsew power bidirectional
rlabel metal5 s -6696 370076 590620 370676 6 vdda1
port 971 nsew power bidirectional
rlabel metal5 s -6696 334076 590620 334676 6 vdda1
port 972 nsew power bidirectional
rlabel metal5 s -6696 298076 590620 298676 6 vdda1
port 973 nsew power bidirectional
rlabel metal5 s -6696 262076 590620 262676 6 vdda1
port 974 nsew power bidirectional
rlabel metal5 s -6696 226076 590620 226676 6 vdda1
port 975 nsew power bidirectional
rlabel metal5 s -6696 190076 590620 190676 6 vdda1
port 976 nsew power bidirectional
rlabel metal5 s -6696 154076 590620 154676 6 vdda1
port 977 nsew power bidirectional
rlabel metal5 s -6696 118076 590620 118676 6 vdda1
port 978 nsew power bidirectional
rlabel metal5 s -6696 82076 590620 82676 6 vdda1
port 979 nsew power bidirectional
rlabel metal5 s -6696 46076 590620 46676 6 vdda1
port 980 nsew power bidirectional
rlabel metal5 s -6696 10076 590620 10676 6 vdda1
port 981 nsew power bidirectional
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 982 nsew power bidirectional
rlabel metal4 s 590020 -5624 590620 709560 6 vssa1
port 983 nsew ground bidirectional
rlabel metal4 s 567004 -5624 567604 709560 6 vssa1
port 984 nsew ground bidirectional
rlabel metal4 s 531004 -5624 531604 709560 6 vssa1
port 985 nsew ground bidirectional
rlabel metal4 s 495004 613200 495604 709560 6 vssa1
port 986 nsew ground bidirectional
rlabel metal4 s 459004 613200 459604 709560 6 vssa1
port 987 nsew ground bidirectional
rlabel metal4 s 423004 -5624 423604 709560 6 vssa1
port 988 nsew ground bidirectional
rlabel metal4 s 387004 613200 387604 709560 6 vssa1
port 989 nsew ground bidirectional
rlabel metal4 s 351004 613200 351604 709560 6 vssa1
port 990 nsew ground bidirectional
rlabel metal4 s 315004 -5624 315604 709560 6 vssa1
port 991 nsew ground bidirectional
rlabel metal4 s 279004 -5624 279604 709560 6 vssa1
port 992 nsew ground bidirectional
rlabel metal4 s 243004 613200 243604 709560 6 vssa1
port 993 nsew ground bidirectional
rlabel metal4 s 207004 613200 207604 709560 6 vssa1
port 994 nsew ground bidirectional
rlabel metal4 s 171004 -5624 171604 709560 6 vssa1
port 995 nsew ground bidirectional
rlabel metal4 s 135004 -5624 135604 709560 6 vssa1
port 996 nsew ground bidirectional
rlabel metal4 s 99004 613200 99604 709560 6 vssa1
port 997 nsew ground bidirectional
rlabel metal4 s 63004 -5624 63604 709560 6 vssa1
port 998 nsew ground bidirectional
rlabel metal4 s 27004 -5624 27604 709560 6 vssa1
port 999 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1
port 1000 nsew ground bidirectional
rlabel metal4 s 495004 460400 495604 549200 6 vssa1
port 1001 nsew ground bidirectional
rlabel metal4 s 459004 460400 459604 549200 6 vssa1
port 1002 nsew ground bidirectional
rlabel metal4 s 387004 460400 387604 549200 6 vssa1
port 1003 nsew ground bidirectional
rlabel metal4 s 351004 460400 351604 549200 6 vssa1
port 1004 nsew ground bidirectional
rlabel metal4 s 243004 460400 243604 549200 6 vssa1
port 1005 nsew ground bidirectional
rlabel metal4 s 207004 460400 207604 549200 6 vssa1
port 1006 nsew ground bidirectional
rlabel metal4 s 99004 460400 99604 549200 6 vssa1
port 1007 nsew ground bidirectional
rlabel metal4 s 495004 307600 495604 396400 6 vssa1
port 1008 nsew ground bidirectional
rlabel metal4 s 459004 307600 459604 396400 6 vssa1
port 1009 nsew ground bidirectional
rlabel metal4 s 387004 307600 387604 396400 6 vssa1
port 1010 nsew ground bidirectional
rlabel metal4 s 351004 307600 351604 396400 6 vssa1
port 1011 nsew ground bidirectional
rlabel metal4 s 243004 307600 243604 396400 6 vssa1
port 1012 nsew ground bidirectional
rlabel metal4 s 207004 307600 207604 396400 6 vssa1
port 1013 nsew ground bidirectional
rlabel metal4 s 99004 307600 99604 396400 6 vssa1
port 1014 nsew ground bidirectional
rlabel metal4 s 495004 154800 495604 243600 6 vssa1
port 1015 nsew ground bidirectional
rlabel metal4 s 459004 154800 459604 243600 6 vssa1
port 1016 nsew ground bidirectional
rlabel metal4 s 387004 154800 387604 243600 6 vssa1
port 1017 nsew ground bidirectional
rlabel metal4 s 351004 154800 351604 243600 6 vssa1
port 1018 nsew ground bidirectional
rlabel metal4 s 243004 154800 243604 243600 6 vssa1
port 1019 nsew ground bidirectional
rlabel metal4 s 207004 154800 207604 243600 6 vssa1
port 1020 nsew ground bidirectional
rlabel metal4 s 99004 154800 99604 243600 6 vssa1
port 1021 nsew ground bidirectional
rlabel metal4 s 495004 -5624 495604 90800 6 vssa1
port 1022 nsew ground bidirectional
rlabel metal4 s 459004 -5624 459604 90800 6 vssa1
port 1023 nsew ground bidirectional
rlabel metal4 s 387004 -5624 387604 90800 6 vssa1
port 1024 nsew ground bidirectional
rlabel metal4 s 351004 -5624 351604 90800 6 vssa1
port 1025 nsew ground bidirectional
rlabel metal4 s 243004 -5624 243604 90800 6 vssa1
port 1026 nsew ground bidirectional
rlabel metal4 s 207004 -5624 207604 90800 6 vssa1
port 1027 nsew ground bidirectional
rlabel metal4 s 99004 -5624 99604 90800 6 vssa1
port 1028 nsew ground bidirectional
rlabel metal5 s -6696 708960 590620 709560 6 vssa1
port 1029 nsew ground bidirectional
rlabel metal5 s -6696 676076 590620 676676 6 vssa1
port 1030 nsew ground bidirectional
rlabel metal5 s -6696 640076 590620 640676 6 vssa1
port 1031 nsew ground bidirectional
rlabel metal5 s -6696 604076 590620 604676 6 vssa1
port 1032 nsew ground bidirectional
rlabel metal5 s -6696 568076 590620 568676 6 vssa1
port 1033 nsew ground bidirectional
rlabel metal5 s -6696 532076 590620 532676 6 vssa1
port 1034 nsew ground bidirectional
rlabel metal5 s -6696 496076 590620 496676 6 vssa1
port 1035 nsew ground bidirectional
rlabel metal5 s -6696 460076 590620 460676 6 vssa1
port 1036 nsew ground bidirectional
rlabel metal5 s -6696 424076 590620 424676 6 vssa1
port 1037 nsew ground bidirectional
rlabel metal5 s -6696 388076 590620 388676 6 vssa1
port 1038 nsew ground bidirectional
rlabel metal5 s -6696 352076 590620 352676 6 vssa1
port 1039 nsew ground bidirectional
rlabel metal5 s -6696 316076 590620 316676 6 vssa1
port 1040 nsew ground bidirectional
rlabel metal5 s -6696 280076 590620 280676 6 vssa1
port 1041 nsew ground bidirectional
rlabel metal5 s -6696 244076 590620 244676 6 vssa1
port 1042 nsew ground bidirectional
rlabel metal5 s -6696 208076 590620 208676 6 vssa1
port 1043 nsew ground bidirectional
rlabel metal5 s -6696 172076 590620 172676 6 vssa1
port 1044 nsew ground bidirectional
rlabel metal5 s -6696 136076 590620 136676 6 vssa1
port 1045 nsew ground bidirectional
rlabel metal5 s -6696 100076 590620 100676 6 vssa1
port 1046 nsew ground bidirectional
rlabel metal5 s -6696 64076 590620 64676 6 vssa1
port 1047 nsew ground bidirectional
rlabel metal5 s -6696 28076 590620 28676 6 vssa1
port 1048 nsew ground bidirectional
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 1049 nsew ground bidirectional
rlabel metal4 s 552604 -7504 553204 711440 6 vdda2
port 1050 nsew power bidirectional
rlabel metal4 s 516604 613200 517204 711440 6 vdda2
port 1051 nsew power bidirectional
rlabel metal4 s 480604 613200 481204 711440 6 vdda2
port 1052 nsew power bidirectional
rlabel metal4 s 444604 -7504 445204 711440 6 vdda2
port 1053 nsew power bidirectional
rlabel metal4 s 408604 -7504 409204 711440 6 vdda2
port 1054 nsew power bidirectional
rlabel metal4 s 372604 613200 373204 711440 6 vdda2
port 1055 nsew power bidirectional
rlabel metal4 s 336604 613200 337204 711440 6 vdda2
port 1056 nsew power bidirectional
rlabel metal4 s 300604 -7504 301204 711440 6 vdda2
port 1057 nsew power bidirectional
rlabel metal4 s 264604 -7504 265204 711440 6 vdda2
port 1058 nsew power bidirectional
rlabel metal4 s 228604 613200 229204 711440 6 vdda2
port 1059 nsew power bidirectional
rlabel metal4 s 192604 -7504 193204 711440 6 vdda2
port 1060 nsew power bidirectional
rlabel metal4 s 156604 -7504 157204 711440 6 vdda2
port 1061 nsew power bidirectional
rlabel metal4 s 120604 613200 121204 711440 6 vdda2
port 1062 nsew power bidirectional
rlabel metal4 s 84604 613200 85204 711440 6 vdda2
port 1063 nsew power bidirectional
rlabel metal4 s 48604 -7504 49204 711440 6 vdda2
port 1064 nsew power bidirectional
rlabel metal4 s 12604 -7504 13204 711440 6 vdda2
port 1065 nsew power bidirectional
rlabel metal4 s 590960 -6564 591560 710500 6 vdda2
port 1066 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2
port 1067 nsew power bidirectional
rlabel metal4 s 516604 460400 517204 549200 6 vdda2
port 1068 nsew power bidirectional
rlabel metal4 s 480604 460400 481204 549200 6 vdda2
port 1069 nsew power bidirectional
rlabel metal4 s 372604 460400 373204 549200 6 vdda2
port 1070 nsew power bidirectional
rlabel metal4 s 336604 460400 337204 549200 6 vdda2
port 1071 nsew power bidirectional
rlabel metal4 s 228604 460400 229204 549200 6 vdda2
port 1072 nsew power bidirectional
rlabel metal4 s 120604 460400 121204 549200 6 vdda2
port 1073 nsew power bidirectional
rlabel metal4 s 84604 460400 85204 549200 6 vdda2
port 1074 nsew power bidirectional
rlabel metal4 s 516604 307600 517204 396400 6 vdda2
port 1075 nsew power bidirectional
rlabel metal4 s 480604 307600 481204 396400 6 vdda2
port 1076 nsew power bidirectional
rlabel metal4 s 372604 307600 373204 396400 6 vdda2
port 1077 nsew power bidirectional
rlabel metal4 s 336604 307600 337204 396400 6 vdda2
port 1078 nsew power bidirectional
rlabel metal4 s 228604 307600 229204 396400 6 vdda2
port 1079 nsew power bidirectional
rlabel metal4 s 120604 307600 121204 396400 6 vdda2
port 1080 nsew power bidirectional
rlabel metal4 s 84604 307600 85204 396400 6 vdda2
port 1081 nsew power bidirectional
rlabel metal4 s 516604 154800 517204 243600 6 vdda2
port 1082 nsew power bidirectional
rlabel metal4 s 480604 154800 481204 243600 6 vdda2
port 1083 nsew power bidirectional
rlabel metal4 s 372604 154800 373204 243600 6 vdda2
port 1084 nsew power bidirectional
rlabel metal4 s 336604 154800 337204 243600 6 vdda2
port 1085 nsew power bidirectional
rlabel metal4 s 228604 154800 229204 243600 6 vdda2
port 1086 nsew power bidirectional
rlabel metal4 s 120604 154800 121204 243600 6 vdda2
port 1087 nsew power bidirectional
rlabel metal4 s 84604 154800 85204 243600 6 vdda2
port 1088 nsew power bidirectional
rlabel metal4 s 516604 -7504 517204 90800 6 vdda2
port 1089 nsew power bidirectional
rlabel metal4 s 480604 -7504 481204 90800 6 vdda2
port 1090 nsew power bidirectional
rlabel metal4 s 372604 -7504 373204 90800 6 vdda2
port 1091 nsew power bidirectional
rlabel metal4 s 336604 -7504 337204 90800 6 vdda2
port 1092 nsew power bidirectional
rlabel metal4 s 228604 -7504 229204 90800 6 vdda2
port 1093 nsew power bidirectional
rlabel metal4 s 120604 -7504 121204 90800 6 vdda2
port 1094 nsew power bidirectional
rlabel metal4 s 84604 -7504 85204 90800 6 vdda2
port 1095 nsew power bidirectional
rlabel metal5 s -7636 709900 591560 710500 6 vdda2
port 1096 nsew power bidirectional
rlabel metal5 s -8576 697676 592500 698276 6 vdda2
port 1097 nsew power bidirectional
rlabel metal5 s -8576 661676 592500 662276 6 vdda2
port 1098 nsew power bidirectional
rlabel metal5 s -8576 625676 592500 626276 6 vdda2
port 1099 nsew power bidirectional
rlabel metal5 s -8576 589676 592500 590276 6 vdda2
port 1100 nsew power bidirectional
rlabel metal5 s -8576 553676 592500 554276 6 vdda2
port 1101 nsew power bidirectional
rlabel metal5 s -8576 517676 592500 518276 6 vdda2
port 1102 nsew power bidirectional
rlabel metal5 s -8576 481676 592500 482276 6 vdda2
port 1103 nsew power bidirectional
rlabel metal5 s -8576 445676 592500 446276 6 vdda2
port 1104 nsew power bidirectional
rlabel metal5 s -8576 409676 592500 410276 6 vdda2
port 1105 nsew power bidirectional
rlabel metal5 s -8576 373676 592500 374276 6 vdda2
port 1106 nsew power bidirectional
rlabel metal5 s -8576 337676 592500 338276 6 vdda2
port 1107 nsew power bidirectional
rlabel metal5 s -8576 301676 592500 302276 6 vdda2
port 1108 nsew power bidirectional
rlabel metal5 s -8576 265676 592500 266276 6 vdda2
port 1109 nsew power bidirectional
rlabel metal5 s -8576 229676 592500 230276 6 vdda2
port 1110 nsew power bidirectional
rlabel metal5 s -8576 193676 592500 194276 6 vdda2
port 1111 nsew power bidirectional
rlabel metal5 s -8576 157676 592500 158276 6 vdda2
port 1112 nsew power bidirectional
rlabel metal5 s -8576 121676 592500 122276 6 vdda2
port 1113 nsew power bidirectional
rlabel metal5 s -8576 85676 592500 86276 6 vdda2
port 1114 nsew power bidirectional
rlabel metal5 s -8576 49676 592500 50276 6 vdda2
port 1115 nsew power bidirectional
rlabel metal5 s -8576 13676 592500 14276 6 vdda2
port 1116 nsew power bidirectional
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 1117 nsew power bidirectional
rlabel metal4 s 591900 -7504 592500 711440 6 vssa2
port 1118 nsew ground bidirectional
rlabel metal4 s 570604 -7504 571204 711440 6 vssa2
port 1119 nsew ground bidirectional
rlabel metal4 s 534604 -7504 535204 711440 6 vssa2
port 1120 nsew ground bidirectional
rlabel metal4 s 498604 613200 499204 711440 6 vssa2
port 1121 nsew ground bidirectional
rlabel metal4 s 462604 613200 463204 711440 6 vssa2
port 1122 nsew ground bidirectional
rlabel metal4 s 426604 -7504 427204 711440 6 vssa2
port 1123 nsew ground bidirectional
rlabel metal4 s 390604 -7504 391204 711440 6 vssa2
port 1124 nsew ground bidirectional
rlabel metal4 s 354604 613200 355204 711440 6 vssa2
port 1125 nsew ground bidirectional
rlabel metal4 s 318604 -7504 319204 711440 6 vssa2
port 1126 nsew ground bidirectional
rlabel metal4 s 282604 -7504 283204 711440 6 vssa2
port 1127 nsew ground bidirectional
rlabel metal4 s 246604 613200 247204 711440 6 vssa2
port 1128 nsew ground bidirectional
rlabel metal4 s 210604 613200 211204 711440 6 vssa2
port 1129 nsew ground bidirectional
rlabel metal4 s 174604 -7504 175204 711440 6 vssa2
port 1130 nsew ground bidirectional
rlabel metal4 s 138604 -7504 139204 711440 6 vssa2
port 1131 nsew ground bidirectional
rlabel metal4 s 102604 613200 103204 711440 6 vssa2
port 1132 nsew ground bidirectional
rlabel metal4 s 66604 613200 67204 711440 6 vssa2
port 1133 nsew ground bidirectional
rlabel metal4 s 30604 -7504 31204 711440 6 vssa2
port 1134 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2
port 1135 nsew ground bidirectional
rlabel metal4 s 498604 460400 499204 549200 6 vssa2
port 1136 nsew ground bidirectional
rlabel metal4 s 462604 460400 463204 549200 6 vssa2
port 1137 nsew ground bidirectional
rlabel metal4 s 354604 460400 355204 549200 6 vssa2
port 1138 nsew ground bidirectional
rlabel metal4 s 246604 460400 247204 549200 6 vssa2
port 1139 nsew ground bidirectional
rlabel metal4 s 210604 460400 211204 549200 6 vssa2
port 1140 nsew ground bidirectional
rlabel metal4 s 102604 460400 103204 549200 6 vssa2
port 1141 nsew ground bidirectional
rlabel metal4 s 66604 460400 67204 549200 6 vssa2
port 1142 nsew ground bidirectional
rlabel metal4 s 498604 307600 499204 396400 6 vssa2
port 1143 nsew ground bidirectional
rlabel metal4 s 462604 307600 463204 396400 6 vssa2
port 1144 nsew ground bidirectional
rlabel metal4 s 354604 307600 355204 396400 6 vssa2
port 1145 nsew ground bidirectional
rlabel metal4 s 246604 307600 247204 396400 6 vssa2
port 1146 nsew ground bidirectional
rlabel metal4 s 210604 307600 211204 396400 6 vssa2
port 1147 nsew ground bidirectional
rlabel metal4 s 102604 307600 103204 396400 6 vssa2
port 1148 nsew ground bidirectional
rlabel metal4 s 66604 307600 67204 396400 6 vssa2
port 1149 nsew ground bidirectional
rlabel metal4 s 498604 154800 499204 243600 6 vssa2
port 1150 nsew ground bidirectional
rlabel metal4 s 462604 154800 463204 243600 6 vssa2
port 1151 nsew ground bidirectional
rlabel metal4 s 354604 154800 355204 243600 6 vssa2
port 1152 nsew ground bidirectional
rlabel metal4 s 246604 154800 247204 243600 6 vssa2
port 1153 nsew ground bidirectional
rlabel metal4 s 210604 154800 211204 243600 6 vssa2
port 1154 nsew ground bidirectional
rlabel metal4 s 102604 154800 103204 243600 6 vssa2
port 1155 nsew ground bidirectional
rlabel metal4 s 66604 154800 67204 243600 6 vssa2
port 1156 nsew ground bidirectional
rlabel metal4 s 498604 -7504 499204 90800 6 vssa2
port 1157 nsew ground bidirectional
rlabel metal4 s 462604 -7504 463204 90800 6 vssa2
port 1158 nsew ground bidirectional
rlabel metal4 s 354604 -7504 355204 90800 6 vssa2
port 1159 nsew ground bidirectional
rlabel metal4 s 246604 -7504 247204 90800 6 vssa2
port 1160 nsew ground bidirectional
rlabel metal4 s 210604 -7504 211204 90800 6 vssa2
port 1161 nsew ground bidirectional
rlabel metal4 s 102604 -7504 103204 90800 6 vssa2
port 1162 nsew ground bidirectional
rlabel metal4 s 66604 -7504 67204 90800 6 vssa2
port 1163 nsew ground bidirectional
rlabel metal5 s -8576 710840 592500 711440 6 vssa2
port 1164 nsew ground bidirectional
rlabel metal5 s -8576 679676 592500 680276 6 vssa2
port 1165 nsew ground bidirectional
rlabel metal5 s -8576 643676 592500 644276 6 vssa2
port 1166 nsew ground bidirectional
rlabel metal5 s -8576 607676 592500 608276 6 vssa2
port 1167 nsew ground bidirectional
rlabel metal5 s -8576 571676 592500 572276 6 vssa2
port 1168 nsew ground bidirectional
rlabel metal5 s -8576 535676 592500 536276 6 vssa2
port 1169 nsew ground bidirectional
rlabel metal5 s -8576 499676 592500 500276 6 vssa2
port 1170 nsew ground bidirectional
rlabel metal5 s -8576 463676 592500 464276 6 vssa2
port 1171 nsew ground bidirectional
rlabel metal5 s -8576 427676 592500 428276 6 vssa2
port 1172 nsew ground bidirectional
rlabel metal5 s -8576 391676 592500 392276 6 vssa2
port 1173 nsew ground bidirectional
rlabel metal5 s -8576 355676 592500 356276 6 vssa2
port 1174 nsew ground bidirectional
rlabel metal5 s -8576 319676 592500 320276 6 vssa2
port 1175 nsew ground bidirectional
rlabel metal5 s -8576 283676 592500 284276 6 vssa2
port 1176 nsew ground bidirectional
rlabel metal5 s -8576 247676 592500 248276 6 vssa2
port 1177 nsew ground bidirectional
rlabel metal5 s -8576 211676 592500 212276 6 vssa2
port 1178 nsew ground bidirectional
rlabel metal5 s -8576 175676 592500 176276 6 vssa2
port 1179 nsew ground bidirectional
rlabel metal5 s -8576 139676 592500 140276 6 vssa2
port 1180 nsew ground bidirectional
rlabel metal5 s -8576 103676 592500 104276 6 vssa2
port 1181 nsew ground bidirectional
rlabel metal5 s -8576 67676 592500 68276 6 vssa2
port 1182 nsew ground bidirectional
rlabel metal5 s -8576 31676 592500 32276 6 vssa2
port 1183 nsew ground bidirectional
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 1184 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 584000 704000
string LEFview TRUE
string GDS_FILE /project/openlane/user_project_wrapper/runs/user_project_wrapper/results/magic/user_project_wrapper.gds
string GDS_END 40528462
string GDS_START 3294246
<< end >>

